
module inverter (di, clk, rstn, do);
 input [15:0] di;
 input clk;
 input rstn;
 output [15:0] do;
  wire \net_Buf-pad-di[15]_IN_to_RIGHT_I326_54_0 ;
  wire \net_Buf-pad-di[15]_RIGHT_LLH11_to_LLH026_27_0 ;
  wire \net_Buf-pad-di[15]_H6W1_to_H6E126_21_0 ;
  wire \net_Buf-pad-di[15]_V6N2_to_V6S220_21_0 ;
  wire \net_Buf-pad-di[15]_V6N2_to_V6S213_21_0 ;
  wire \net_Buf-pad-di[15]_N13_to_S1312_21_0 ;
  wire \net_Buf-pad-di[15]_S0_F_B1_to_F112_21_0 ;
  wire net_VCC_X_to_S0_X7_21_0;
  wire net_VCC_V6S1_to_V6N113_21_0;
  wire net_VCC_N7_to_S712_21_0;
  wire net_VCC_S0_F_B2_to_F212_21_0;
  wire net_VCC_S0_G_B2_to_G212_21_0;
  wire net_VCC_V6S2_to_V6M210_21_0;
  wire net_VCC_S16_to_N1611_21_0;
  wire net_VCC_S0_F_B2_to_F211_21_0;
  wire net_VCC_S0_G_B2_to_G211_21_0;
  wire net_VCC_N14_to_S146_21_0;
  wire net_VCC_N14_to_S145_21_0;
  wire net_VCC_S1_F_B2_to_F25_21_0;
  wire net_VCC_S1_G_B2_to_G25_21_0;
  wire net_VCC_S13_to_N138_21_0;
  wire net_VCC_S1_F_B2_to_F28_21_0;
  wire net_VCC_S1_G_B2_to_G28_21_0;
  wire net_VCC_S13_to_N139_21_0;
  wire net_VCC_S1_F_B2_to_F29_21_0;
  wire net_VCC_S1_G_B2_to_G29_21_0;
  wire net_VCC_N1_to_S16_21_0;
  wire net_VCC_N1_to_S15_21_0;
  wire net_VCC_S0_F_B2_to_F25_21_0;
  wire net_VCC_S0_G_B2_to_G25_21_0;
  wire net_VCC_V6N7_to_V6M74_21_0;
  wire net_VCC_S0_F_B2_to_F24_21_0;
  wire net_VCC_S0_G_B2_to_G24_21_0;
  wire net_VCC_S0_F_B2_to_F26_21_0;
  wire net_VCC_S0_G_B2_to_G26_21_0;
  wire \net_Buf-pad-di[14]_IN_to_TOP_I11_21_0 ;
  wire \net_Buf-pad-di[14]_TOP_V6C2_to_V6N25_21_0 ;
  wire \net_Buf-pad-di[14]_V6S2_to_V6N211_21_0 ;
  wire \net_Buf-pad-di[14]_S14_to_N1412_21_0 ;
  wire \net_Buf-pad-di[14]_S0_G_B1_to_G112_21_0 ;
  wire \net_Buf-pad-di[13]_IN_to_TOP_I11_35_0 ;
  wire \net_Buf-pad-di[13]_TOP_H6W0_to_TOP_H6E01_29_0 ;
  wire \net_Buf-pad-di[13]_TOP_H6W0_to_TOP_H6E01_22_0 ;
  wire \net_Buf-pad-di[13]_TOP_V6D8_to_V6N86_22_0 ;
  wire \net_Buf-pad-di[13]_V6S8_to_V6N812_22_0 ;
  wire \net_Buf-pad-di[13]_W8_to_E812_21_0 ;
  wire \net_Buf-pad-di[13]_N12_to_S1211_21_0 ;
  wire \net_Buf-pad-di[13]_S0_F_B1_to_F111_21_0 ;
  wire \net_Buf-pad-di[12]_IN_to_TOP_I21_40_0 ;
  wire \net_Buf-pad-di[12]_TOP_H6W3_to_TOP_H6E31_34_0 ;
  wire \net_Buf-pad-di[12]_TOP_H6W3_to_TOP_H6E31_27_0 ;
  wire \net_Buf-pad-di[12]_TOP_V6S2_to_V6M24_27_0 ;
  wire \net_Buf-pad-di[12]_H6W2_to_H6E24_21_0 ;
  wire \net_Buf-pad-di[12]_V6S3_to_V6N310_21_0 ;
  wire \net_Buf-pad-di[12]_S22_to_N2211_21_0 ;
  wire \net_Buf-pad-di[12]_S0_G_B1_to_G111_21_0 ;
  wire \net_Buf-pad-di[11]_IN_to_TOP_I11_40_0 ;
  wire \net_Buf-pad-di[11]_TOP_H6W2_to_TOP_H6E21_34_0 ;
  wire \net_Buf-pad-di[11]_TOP_H6W2_to_TOP_H6E21_27_0 ;
  wire \net_Buf-pad-di[11]_TOP_V6D4_to_V6N46_27_0 ;
  wire \net_Buf-pad-di[11]_H6W8_to_H6E86_21_0 ;
  wire \net_Buf-pad-di[11]_N9_to_S95_21_0 ;
  wire \net_Buf-pad-di[11]_S1_F_B1_to_F15_21_0 ;
  wire \net_Buf-pad-di[10]_IN_to_TOP_I21_42_0 ;
  wire \net_Buf-pad-di[10]_TOP_LLH6_to_TOP_LLH01_22_0 ;
  wire \net_Buf-pad-di[10]_TOP_H6W4_to_TOP_H6C41_20_0 ;
  wire \net_Buf-pad-di[10]_TOP_LLV8_to_LLV05_20_0 ;
  wire \net_Buf-pad-di[10]_E9_to_W95_21_0 ;
  wire \net_Buf-pad-di[10]_S1_G_B1_to_G15_21_0 ;
  wire \net_Buf-pad-di[9]_IN_to_TOP_I11_44_0 ;
  wire \net_Buf-pad-di[9]_TOP_LLH0_to_TOP_LLH61_24_0 ;
  wire \net_Buf-pad-di[9]_TOP_H6W3_to_TOP_H6M31_21_0 ;
  wire \net_Buf-pad-di[9]_TOP_V6S8_to_V6N87_21_0 ;
  wire \net_Buf-pad-di[9]_S5_to_N58_21_0 ;
  wire \net_Buf-pad-di[9]_S1_F_B1_to_F18_21_0 ;
  wire \net_Buf-pad-di[8]_IN_to_TOP_I21_47_0 ;
  wire \net_Buf-pad-di[8]_TOP_H6W3_to_TOP_H6E31_40_0 ;
  wire \net_Buf-pad-di[8]_TOP_V6S10_to_V6N107_40_0 ;
  wire \net_Buf-pad-di[8]_H6W4_to_H6E47_34_0 ;
  wire \net_Buf-pad-di[8]_H6W4_to_H6E47_27_0 ;
  wire \net_Buf-pad-di[8]_H6W4_to_H6E47_21_0 ;
  wire \net_Buf-pad-di[8]_S3_to_N38_21_0 ;
  wire \net_Buf-pad-di[8]_S1_G_B1_to_G18_21_0 ;
  wire \net_Buf-pad-di[7]_IN_to_TOP_I11_47_0 ;
  wire \net_Buf-pad-di[7]_TOP_H6W1_to_TOP_H6E11_40_0 ;
  wire \net_Buf-pad-di[7]_TOP_H6W1_to_TOP_H6E11_34_0 ;
  wire \net_Buf-pad-di[7]_TOP_H6W1_to_TOP_H6E11_27_0 ;
  wire \net_Buf-pad-di[7]_TOP_V6D6_to_V6N66_27_0 ;
  wire \net_Buf-pad-di[7]_H6W10_to_H6E106_21_0 ;
  wire \net_Buf-pad-di[7]_V6S10_to_V6M109_21_0 ;
  wire \net_Buf-pad-di[7]_S1_F_B1_to_F19_21_0 ;
  wire \net_Buf-pad-di[6]_IN_to_TOP_I21_48_0 ;
  wire \net_Buf-pad-di[6]_TOP_LLH6_to_TOP_LLH61_22_0 ;
  wire \net_Buf-pad-di[6]_TOP_V6S6_to_V6N67_22_0 ;
  wire \net_Buf-pad-di[6]_V6S6_to_V6M610_22_0 ;
  wire \net_Buf-pad-di[6]_W14_to_E1410_21_0 ;
  wire \net_Buf-pad-di[6]_N18_to_S189_21_0 ;
  wire \net_Buf-pad-di[6]_S1_G_B1_to_G19_21_0 ;
  wire \net_Buf-pad-di[5]_IN_to_TOP_I11_50_0 ;
  wire \net_Buf-pad-di[5]_TOP_LLH0_to_TOP_LLH61_18_0 ;
  wire \net_Buf-pad-di[5]_TOP_H6E2_to_TOP_H6M21_21_0 ;
  wire \net_Buf-pad-di[5]_TOP_V6D10_to_V6N106_21_0 ;
  wire \net_Buf-pad-di[5]_N17_to_S175_21_0 ;
  wire \net_Buf-pad-di[5]_S0_F_B1_to_F15_21_0 ;
  wire \net_Buf-pad-di[4]_IN_to_TOP_I21_53_0 ;
  wire \net_Buf-pad-di[4]_TOP_LLH0_to_TOP_LLH61_21_0 ;
  wire \net_Buf-pad-di[4]_TOP_V6D8_to_V6N86_21_0 ;
  wire \net_Buf-pad-di[4]_N5_to_S55_21_0 ;
  wire \net_Buf-pad-di[4]_S0_G_B1_to_G15_21_0 ;
  wire \net_Buf-pad-di[3]_IN_to_TOP_I11_53_0 ;
  wire \net_Buf-pad-di[3]_TOP_LLH6_to_TOP_LLH01_21_0 ;
  wire \net_Buf-pad-di[3]_TOP_V6S6_to_V6M64_21_0 ;
  wire \net_Buf-pad-di[3]_S0_F_B1_to_F14_21_0 ;
  wire \net_Buf-pad-di[2]_IN_to_RIGHT_I14_54_0 ;
  wire \net_Buf-pad-di[2]_RIGHT_LLH4_to_LLH04_20_0 ;
  wire \net_Buf-pad-di[2]_E22_to_W224_21_0 ;
  wire \net_Buf-pad-di[2]_S0_G_B1_to_G14_21_0 ;
  wire \net_Buf-pad-di[1]_IN_to_RIGHT_I16_54_0 ;
  wire \net_Buf-pad-di[1]_RIGHT_LLH4_to_LLH06_20_0 ;
  wire \net_Buf-pad-di[1]_E22_to_W226_21_0 ;
  wire \net_Buf-pad-di[1]_S0_F_B1_to_F16_21_0 ;
  wire \net_Buf-pad-di[0]_IN_to_RIGHT_I18_54_0 ;
  wire \net_Buf-pad-di[0]_RIGHT_LLH4_to_LLH08_20_0 ;
  wire \net_Buf-pad-di[0]_V6N0_to_V6M05_20_0 ;
  wire \net_Buf-pad-di[0]_E1_to_W15_21_0 ;
  wire \net_Buf-pad-di[0]_S23_to_N236_21_0 ;
  wire \net_Buf-pad-di[0]_S0_G_B1_to_G16_21_0 ;
  wire \net_Buf-pad-clk_GCLKOUT_to_CLKB_CLKPAD135_28_0 ;
  wire \net_Buf-pad-clk_CLKB_GCLKBUF1_IN_to_IN35_28_0 ;
  wire \net_do_reg[15]_XQ_to_S0_XQ12_21_0 ;
  wire \net_do_reg[15]_LLH6_to_LLH612_8_0 ;
  wire \net_do_reg[15]_H6W3_to_LEFT_H6E312_2_0 ;
  wire \net_do_reg[15]_LEFT_V6S3_to_LEFT_V6N319_2_0 ;
  wire \net_do_reg[15]_LEFT_E20_to_W2019_3_0 ;
  wire \net_do_reg[15]_N19_to_S1917_3_0 ;
  wire \net_do_reg[15]_W21_to_LEFT_E2117_2_0 ;
  wire \net_do_reg[15]_LEFT_O2_to_OUT17_2_0 ;
  wire \net_do_reg[14]_YQ_to_S0_YQ12_21_0 ;
  wire \net_do_reg[14]_LLH0_to_LLH012_8_0 ;
  wire \net_do_reg[14]_H6W0_to_LEFT_H6E012_2_0 ;
  wire \net_do_reg[14]_LEFT_V6S0_to_LEFT_V6M015_2_0 ;
  wire \net_do_reg[14]_LEFT_E1_to_W115_3_0 ;
  wire \net_do_reg[14]_N20_to_S2014_3_0 ;
  wire \net_do_reg[14]_W22_to_LEFT_E2214_2_0 ;
  wire \net_do_reg[14]_LEFT_O2_to_OUT14_2_0 ;
  wire \net_do_reg[13]_XQ_to_S0_XQ11_21_0 ;
  wire \net_do_reg[13]_LLH6_to_LEFT_LLH011_2_0 ;
  wire \net_do_reg[13]_LEFT_V6S0_to_LEFT_V6N017_2_0 ;
  wire \net_do_reg[13]_LEFT_E2_to_W217_3_0 ;
  wire \net_do_reg[13]_N1_to_S116_3_0 ;
  wire \net_do_reg[13]_W7_to_LEFT_E716_2_0 ;
  wire \net_do_reg[13]_LEFT_O1_to_OUT16_2_0 ;
  wire \net_do_reg[12]_YQ_to_S0_YQ11_21_0 ;
  wire \net_do_reg[12]_LLH0_to_LEFT_LLH611_2_0 ;
  wire \net_do_reg[12]_LEFT_V6S3_to_LEFT_V6M314_2_0 ;
  wire \net_do_reg[12]_LEFT_E19_to_W1914_3_0 ;
  wire \net_do_reg[12]_N14_to_S1413_3_0 ;
  wire \net_do_reg[12]_W12_to_LEFT_E1213_2_0 ;
  wire \net_do_reg[12]_LEFT_O2_to_OUT13_2_0 ;
  wire \net_do_reg[11]_XQ_to_S1_XQ5_21_0 ;
  wire \net_do_reg[11]_H6W2_to_H6E25_14_0 ;
  wire \net_do_reg[11]_H6W2_to_H6E25_8_0 ;
  wire \net_do_reg[11]_H6W2_to_LEFT_H6E25_2_0 ;
  wire \net_do_reg[11]_LEFT_V6S2_to_LEFT_V6N211_2_0 ;
  wire \net_do_reg[11]_LEFT_V6S2_to_LEFT_V6M214_2_0 ;
  wire \net_do_reg[11]_LEFT_E16_to_W1614_3_0 ;
  wire \net_do_reg[11]_N15_to_S1513_3_0 ;
  wire \net_do_reg[11]_W17_to_LEFT_E1713_2_0 ;
  wire \net_do_reg[11]_LEFT_O3_to_OUT13_2_0 ;
  wire \net_do_reg[10]_YQ_to_S1_YQ5_21_0 ;
  wire \net_do_reg[10]_H6W3_to_H6E35_14_0 ;
  wire \net_do_reg[10]_V6S0_to_V6N011_14_0 ;
  wire \net_do_reg[10]_H6W0_to_H6E011_8_0 ;
  wire \net_do_reg[10]_V6S1_to_V6M114_8_0 ;
  wire \net_do_reg[10]_H6W1_to_LEFT_H6E114_2_0 ;
  wire \net_do_reg[10]_LEFT_O1_to_OUT14_2_0 ;
  wire \net_do_reg[9]_XQ_to_S1_XQ8_21_0 ;
  wire \net_do_reg[9]_LLH6_to_LLH68_8_0 ;
  wire \net_do_reg[9]_H6W2_to_LEFT_H6E28_2_0 ;
  wire \net_do_reg[9]_LEFT_E12_to_W128_3_0 ;
  wire \net_do_reg[9]_S14_to_N149_3_0 ;
  wire \net_do_reg[9]_W19_to_LEFT_E199_2_0 ;
  wire \net_do_reg[9]_LEFT_O2_to_OUT9_2_0 ;
  wire \net_do_reg[8]_YQ_to_S1_YQ8_21_0 ;
  wire \net_do_reg[8]_LLH0_to_LLH08_8_0 ;
  wire \net_do_reg[8]_H6W0_to_LEFT_H6E08_2_0 ;
  wire \net_do_reg[8]_LEFT_E3_to_W38_3_0 ;
  wire \net_do_reg[8]_S21_to_N219_3_0 ;
  wire \net_do_reg[8]_W22_to_LEFT_E229_2_0 ;
  wire \net_do_reg[8]_LEFT_O3_to_OUT9_2_0 ;
  wire \net_do_reg[7]_XQ_to_S1_XQ9_21_0 ;
  wire \net_do_reg[7]_LLH6_to_LEFT_LLH09_2_0 ;
  wire \net_do_reg[7]_LEFT_E0_to_W09_3_0 ;
  wire \net_do_reg[7]_S2_to_N210_3_0 ;
  wire \net_do_reg[7]_W7_to_LEFT_E710_2_0 ;
  wire \net_do_reg[7]_LEFT_O1_to_OUT10_2_0 ;
  wire \net_do_reg[6]_YQ_to_S1_YQ9_21_0 ;
  wire \net_do_reg[6]_LLH0_to_LEFT_LLH69_2_0 ;
  wire \net_do_reg[6]_LEFT_E23_to_W239_3_0 ;
  wire \net_do_reg[6]_S17_to_N1710_3_0 ;
  wire \net_do_reg[6]_W18_to_LEFT_E1810_2_0 ;
  wire \net_do_reg[6]_LEFT_O2_to_OUT10_2_0 ;
  wire \net_do_reg[5]_XQ_to_S0_XQ5_21_0 ;
  wire \net_do_reg[5]_LLH0_to_LLH05_8_0 ;
  wire \net_do_reg[5]_H6W1_to_H6M15_5_0 ;
  wire \net_do_reg[5]_V6S1_to_V6M18_5_0 ;
  wire \net_do_reg[5]_H6W1_to_LEFT_H6M18_2_0 ;
  wire \net_do_reg[5]_LEFT_O1_to_OUT8_2_0 ;
  wire \net_do_reg[4]_YQ_to_S0_YQ5_21_0 ;
  wire \net_do_reg[4]_LLH6_to_LLH65_8_0 ;
  wire \net_do_reg[4]_H6W3_to_LEFT_H6E35_2_0 ;
  wire \net_do_reg[4]_LEFT_V6S3_to_LEFT_V6M38_2_0 ;
  wire \net_do_reg[4]_LEFT_E22_to_W228_3_0 ;
  wire \net_do_reg[4]_S20_to_N209_3_0 ;
  wire \net_do_reg[4]_W1_to_LEFT_E19_2_0 ;
  wire \net_do_reg[4]_LEFT_O1_to_OUT9_2_0 ;
  wire \net_do_reg[3]_XQ_to_S0_XQ4_21_0 ;
  wire \net_do_reg[3]_LLH0_to_LLH04_8_0 ;
  wire \net_do_reg[3]_H6W1_to_LEFT_H6E14_2_0 ;
  wire \net_do_reg[3]_LEFT_O1_to_OUT4_2_0 ;
  wire \net_do_reg[2]_YQ_to_S0_YQ4_21_0 ;
  wire \net_do_reg[2]_LLH6_to_LEFT_LLH04_2_0 ;
  wire \net_do_reg[2]_LEFT_E8_to_W84_3_0 ;
  wire \net_do_reg[2]_S10_to_N105_3_0 ;
  wire \net_do_reg[2]_W15_to_LEFT_E155_2_0 ;
  wire \net_do_reg[2]_LEFT_O3_to_OUT5_2_0 ;
  wire \net_do_reg[1]_XQ_to_S0_XQ6_21_0 ;
  wire \net_do_reg[1]_LLH6_to_LEFT_LLH06_2_0 ;
  wire \net_do_reg[1]_LEFT_O1_to_OUT6_2_0 ;
  wire \net_do_reg[0]_YQ_to_S0_YQ6_21_0 ;
  wire \net_do_reg[0]_LLH0_to_LEFT_LLH66_2_0 ;
  wire \net_do_reg[0]_LEFT_O2_to_OUT6_2_0 ;
  wire \net_IBuf-clkpad-clk_OUT_to_CLKB_GCLK1_PW35_28_0 ;
  wire \net_IBuf-clkpad-clk_CLKB_GCLK1_to_CLKC_GCLK118_28_0 ;
  wire \net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK112_28_0 ;
  wire \net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK112_21_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK12_21_0 ;
  wire \net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK111_21_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK11_21_0 ;
  wire \net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK15_21_0 ;
  wire \net_IBuf-clkpad-clk_S1_CLK_B_to_CLK5_21_0 ;
  wire \net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK18_21_0 ;
  wire \net_IBuf-clkpad-clk_S1_CLK_B_to_CLK8_21_0 ;
  wire \net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK19_21_0 ;
  wire \net_IBuf-clkpad-clk_S1_CLK_B_to_CLK9_21_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK5_21_0 ;
  wire \net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK14_21_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK4_21_0 ;
  wire \net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK16_21_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK6_21_0 ;
  wire \net_Buf-pad-rstn_IN_to_RIGHT_I35_54_0 ;
  wire \net_Buf-pad-rstn_RIGHT_LLH2_to_LLH05_18_0 ;
  wire \net_Buf-pad-rstn_H6E1_to_H6M15_21_0 ;
  wire \net_Buf-pad-rstn_V6S1_to_V6N111_21_0 ;
  wire \net_Buf-pad-rstn_V6S1_to_V6D112_21_0 ;
  wire \net_Buf-pad-rstn_S0_SR_B_to_SR12_21_0 ;
  wire \net_Buf-pad-rstn_S0_SR_B_to_SR11_21_0 ;
  wire \net_Buf-pad-rstn_S1_SR_B_to_SR5_21_0 ;
  wire \net_Buf-pad-rstn_S1_SR_B_to_SR8_21_0 ;
  wire \net_Buf-pad-rstn_S1_SR_B_to_SR9_21_0 ;
  wire \net_Buf-pad-rstn_S0_SR_B_to_SR5_21_0 ;
  wire \net_Buf-pad-rstn_V6N1_to_V6A14_21_0 ;
  wire \net_Buf-pad-rstn_S0_SR_B_to_SR4_21_0 ;
  wire \net_Buf-pad-rstn_S0_SR_B_to_SR6_21_0 ;


  defparam iSlice__0___inst.ckinv.CONF = "1";
  defparam iSlice__0___inst.dxmux.CONF = "1";
  defparam iSlice__0___inst.dymux.CONF = "1";
  defparam iSlice__0___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__0___inst.ffx.TYPE = "#FF";
  defparam iSlice__0___inst.ffy.TYPE = "#FF";
  defparam iSlice__0___inst.fxmux.CONF = "F";
  defparam iSlice__0___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__0___inst.gymux.CONF = "G";
  defparam iSlice__0___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__0___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__0___inst.srffmux.CONF = "0";
  defparam iSlice__0___inst.srmux.CONF = "SR_B";
  defparam iSlice__0___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__0___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__0___inst.f.INIT = 16'h5;
  defparam iSlice__0___inst.g.INIT = 16'h5;
  SLICE iSlice__0___inst (
    .CIN(),
    .SR(\net_Buf-pad-rstn_S0_SR_B_to_SR12_21_0 ),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK12_21_0 ),
    .CE(),
    .BX(),
    .F1(\net_Buf-pad-di[15]_S0_F_B1_to_F112_21_0 ),
    .F2(net_VCC_S0_F_B2_to_F212_21_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-di[14]_S0_G_B1_to_G112_21_0 ),
    .G2(net_VCC_S0_G_B2_to_G212_21_0),
    .G3(),
    .G4(),
    .XQ(\net_do_reg[15]_XQ_to_S0_XQ12_21_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_do_reg[14]_YQ_to_S0_YQ12_21_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__1___inst.ckinv.CONF = "1";
  defparam iSlice__1___inst.dxmux.CONF = "1";
  defparam iSlice__1___inst.dymux.CONF = "1";
  defparam iSlice__1___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__1___inst.ffx.TYPE = "#FF";
  defparam iSlice__1___inst.ffy.TYPE = "#FF";
  defparam iSlice__1___inst.fxmux.CONF = "F";
  defparam iSlice__1___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__1___inst.gymux.CONF = "G";
  defparam iSlice__1___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__1___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__1___inst.srffmux.CONF = "0";
  defparam iSlice__1___inst.srmux.CONF = "SR_B";
  defparam iSlice__1___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__1___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__1___inst.f.INIT = 16'h5;
  defparam iSlice__1___inst.g.INIT = 16'h5;
  SLICE iSlice__1___inst (
    .CIN(),
    .SR(\net_Buf-pad-rstn_S0_SR_B_to_SR11_21_0 ),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK11_21_0 ),
    .CE(),
    .BX(),
    .F1(\net_Buf-pad-di[13]_S0_F_B1_to_F111_21_0 ),
    .F2(net_VCC_S0_F_B2_to_F211_21_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-di[12]_S0_G_B1_to_G111_21_0 ),
    .G2(net_VCC_S0_G_B2_to_G211_21_0),
    .G3(),
    .G4(),
    .XQ(\net_do_reg[13]_XQ_to_S0_XQ11_21_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_do_reg[12]_YQ_to_S0_YQ11_21_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__2___inst.ckinv.CONF = "1";
  defparam iSlice__2___inst.dxmux.CONF = "1";
  defparam iSlice__2___inst.dymux.CONF = "1";
  defparam iSlice__2___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__2___inst.ffx.TYPE = "#FF";
  defparam iSlice__2___inst.ffy.TYPE = "#FF";
  defparam iSlice__2___inst.fxmux.CONF = "F";
  defparam iSlice__2___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__2___inst.gymux.CONF = "G";
  defparam iSlice__2___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__2___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__2___inst.srffmux.CONF = "0";
  defparam iSlice__2___inst.srmux.CONF = "SR_B";
  defparam iSlice__2___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__2___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__2___inst.f.INIT = 16'h5;
  defparam iSlice__2___inst.g.INIT = 16'h5;
  SLICE iSlice__2___inst (
    .CIN(),
    .SR(\net_Buf-pad-rstn_S1_SR_B_to_SR5_21_0 ),
    .CLK(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK5_21_0 ),
    .CE(),
    .BX(),
    .F1(\net_Buf-pad-di[11]_S1_F_B1_to_F15_21_0 ),
    .F2(net_VCC_S1_F_B2_to_F25_21_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-di[10]_S1_G_B1_to_G15_21_0 ),
    .G2(net_VCC_S1_G_B2_to_G25_21_0),
    .G3(),
    .G4(),
    .XQ(\net_do_reg[11]_XQ_to_S1_XQ5_21_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_do_reg[10]_YQ_to_S1_YQ5_21_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__3___inst.ckinv.CONF = "1";
  defparam iSlice__3___inst.dxmux.CONF = "1";
  defparam iSlice__3___inst.dymux.CONF = "1";
  defparam iSlice__3___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__3___inst.ffx.TYPE = "#FF";
  defparam iSlice__3___inst.ffy.TYPE = "#FF";
  defparam iSlice__3___inst.fxmux.CONF = "F";
  defparam iSlice__3___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__3___inst.gymux.CONF = "G";
  defparam iSlice__3___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__3___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__3___inst.srffmux.CONF = "0";
  defparam iSlice__3___inst.srmux.CONF = "SR_B";
  defparam iSlice__3___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__3___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__3___inst.f.INIT = 16'h5;
  defparam iSlice__3___inst.g.INIT = 16'h5;
  SLICE iSlice__3___inst (
    .CIN(),
    .SR(\net_Buf-pad-rstn_S1_SR_B_to_SR8_21_0 ),
    .CLK(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK8_21_0 ),
    .CE(),
    .BX(),
    .F1(\net_Buf-pad-di[9]_S1_F_B1_to_F18_21_0 ),
    .F2(net_VCC_S1_F_B2_to_F28_21_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-di[8]_S1_G_B1_to_G18_21_0 ),
    .G2(net_VCC_S1_G_B2_to_G28_21_0),
    .G3(),
    .G4(),
    .XQ(\net_do_reg[9]_XQ_to_S1_XQ8_21_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_do_reg[8]_YQ_to_S1_YQ8_21_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__4___inst.ckinv.CONF = "1";
  defparam iSlice__4___inst.dxmux.CONF = "1";
  defparam iSlice__4___inst.dymux.CONF = "1";
  defparam iSlice__4___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__4___inst.ffx.TYPE = "#FF";
  defparam iSlice__4___inst.ffy.TYPE = "#FF";
  defparam iSlice__4___inst.fxmux.CONF = "F";
  defparam iSlice__4___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__4___inst.gymux.CONF = "G";
  defparam iSlice__4___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__4___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__4___inst.srffmux.CONF = "0";
  defparam iSlice__4___inst.srmux.CONF = "SR_B";
  defparam iSlice__4___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__4___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__4___inst.f.INIT = 16'h5;
  defparam iSlice__4___inst.g.INIT = 16'h5;
  SLICE iSlice__4___inst (
    .CIN(),
    .SR(\net_Buf-pad-rstn_S1_SR_B_to_SR9_21_0 ),
    .CLK(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK9_21_0 ),
    .CE(),
    .BX(),
    .F1(\net_Buf-pad-di[7]_S1_F_B1_to_F19_21_0 ),
    .F2(net_VCC_S1_F_B2_to_F29_21_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-di[6]_S1_G_B1_to_G19_21_0 ),
    .G2(net_VCC_S1_G_B2_to_G29_21_0),
    .G3(),
    .G4(),
    .XQ(\net_do_reg[7]_XQ_to_S1_XQ9_21_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_do_reg[6]_YQ_to_S1_YQ9_21_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__5___inst.ckinv.CONF = "1";
  defparam iSlice__5___inst.dxmux.CONF = "1";
  defparam iSlice__5___inst.dymux.CONF = "1";
  defparam iSlice__5___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__5___inst.ffx.TYPE = "#FF";
  defparam iSlice__5___inst.ffy.TYPE = "#FF";
  defparam iSlice__5___inst.fxmux.CONF = "F";
  defparam iSlice__5___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__5___inst.gymux.CONF = "G";
  defparam iSlice__5___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__5___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__5___inst.srffmux.CONF = "0";
  defparam iSlice__5___inst.srmux.CONF = "SR_B";
  defparam iSlice__5___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__5___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__5___inst.f.INIT = 16'h5;
  defparam iSlice__5___inst.g.INIT = 16'h5;
  SLICE iSlice__5___inst (
    .CIN(),
    .SR(\net_Buf-pad-rstn_S0_SR_B_to_SR5_21_0 ),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK5_21_0 ),
    .CE(),
    .BX(),
    .F1(\net_Buf-pad-di[5]_S0_F_B1_to_F15_21_0 ),
    .F2(net_VCC_S0_F_B2_to_F25_21_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-di[4]_S0_G_B1_to_G15_21_0 ),
    .G2(net_VCC_S0_G_B2_to_G25_21_0),
    .G3(),
    .G4(),
    .XQ(\net_do_reg[5]_XQ_to_S0_XQ5_21_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_do_reg[4]_YQ_to_S0_YQ5_21_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__6___inst.ckinv.CONF = "1";
  defparam iSlice__6___inst.dxmux.CONF = "1";
  defparam iSlice__6___inst.dymux.CONF = "1";
  defparam iSlice__6___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__6___inst.ffx.TYPE = "#FF";
  defparam iSlice__6___inst.ffy.TYPE = "#FF";
  defparam iSlice__6___inst.fxmux.CONF = "F";
  defparam iSlice__6___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__6___inst.gymux.CONF = "G";
  defparam iSlice__6___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__6___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__6___inst.srffmux.CONF = "0";
  defparam iSlice__6___inst.srmux.CONF = "SR_B";
  defparam iSlice__6___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__6___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__6___inst.f.INIT = 16'h5;
  defparam iSlice__6___inst.g.INIT = 16'h5;
  SLICE iSlice__6___inst (
    .CIN(),
    .SR(\net_Buf-pad-rstn_S0_SR_B_to_SR4_21_0 ),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK4_21_0 ),
    .CE(),
    .BX(),
    .F1(\net_Buf-pad-di[3]_S0_F_B1_to_F14_21_0 ),
    .F2(net_VCC_S0_F_B2_to_F24_21_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-di[2]_S0_G_B1_to_G14_21_0 ),
    .G2(net_VCC_S0_G_B2_to_G24_21_0),
    .G3(),
    .G4(),
    .XQ(\net_do_reg[3]_XQ_to_S0_XQ4_21_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_do_reg[2]_YQ_to_S0_YQ4_21_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__7___inst.ckinv.CONF = "1";
  defparam iSlice__7___inst.dxmux.CONF = "1";
  defparam iSlice__7___inst.dymux.CONF = "1";
  defparam iSlice__7___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__7___inst.ffx.TYPE = "#FF";
  defparam iSlice__7___inst.ffy.TYPE = "#FF";
  defparam iSlice__7___inst.fxmux.CONF = "F";
  defparam iSlice__7___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__7___inst.gymux.CONF = "G";
  defparam iSlice__7___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__7___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__7___inst.srffmux.CONF = "0";
  defparam iSlice__7___inst.srmux.CONF = "SR_B";
  defparam iSlice__7___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__7___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__7___inst.f.INIT = 16'h5;
  defparam iSlice__7___inst.g.INIT = 16'h5;
  SLICE iSlice__7___inst (
    .CIN(),
    .SR(\net_Buf-pad-rstn_S0_SR_B_to_SR6_21_0 ),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK6_21_0 ),
    .CE(),
    .BX(),
    .F1(\net_Buf-pad-di[1]_S0_F_B1_to_F16_21_0 ),
    .F2(net_VCC_S0_F_B2_to_F26_21_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-di[0]_S0_G_B1_to_G16_21_0 ),
    .G2(net_VCC_S0_G_B2_to_G26_21_0),
    .G3(),
    .G4(),
    .XQ(\net_do_reg[1]_XQ_to_S0_XQ6_21_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_do_reg[0]_YQ_to_S0_YQ6_21_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__8___inst.f.CONF = "#LUT:D=1";
  defparam iSlice__8___inst.fxmux.CONF = "F";
  defparam iSlice__8___inst.xused.CONF = "0";
  defparam iSlice__8___inst.f.INIT = 16'hffff;
  SLICE iSlice__8___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(),
    .F2(),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(net_VCC_X_to_S0_X7_21_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam \di[15]_inst .imux.CONF = "1";
  defparam \di[15]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[15]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[15]_IN_to_RIGHT_I326_54_0 ),
    .IQ(),
    .PAD(di[15])
  );

  defparam \di[14]_inst .imux.CONF = "1";
  defparam \di[14]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[14]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[14]_IN_to_TOP_I11_21_0 ),
    .IQ(),
    .PAD(di[14])
  );

  defparam \di[13]_inst .imux.CONF = "1";
  defparam \di[13]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[13]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[13]_IN_to_TOP_I11_35_0 ),
    .IQ(),
    .PAD(di[13])
  );

  defparam \di[12]_inst .imux.CONF = "1";
  defparam \di[12]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[12]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[12]_IN_to_TOP_I21_40_0 ),
    .IQ(),
    .PAD(di[12])
  );

  defparam \di[11]_inst .imux.CONF = "1";
  defparam \di[11]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[11]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[11]_IN_to_TOP_I11_40_0 ),
    .IQ(),
    .PAD(di[11])
  );

  defparam \di[10]_inst .imux.CONF = "1";
  defparam \di[10]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[10]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[10]_IN_to_TOP_I21_42_0 ),
    .IQ(),
    .PAD(di[10])
  );

  defparam \di[9]_inst .imux.CONF = "1";
  defparam \di[9]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[9]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[9]_IN_to_TOP_I11_44_0 ),
    .IQ(),
    .PAD(di[9])
  );

  defparam \di[8]_inst .imux.CONF = "1";
  defparam \di[8]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[8]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[8]_IN_to_TOP_I21_47_0 ),
    .IQ(),
    .PAD(di[8])
  );

  defparam \di[7]_inst .imux.CONF = "1";
  defparam \di[7]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[7]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[7]_IN_to_TOP_I11_47_0 ),
    .IQ(),
    .PAD(di[7])
  );

  defparam \di[6]_inst .imux.CONF = "1";
  defparam \di[6]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[6]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[6]_IN_to_TOP_I21_48_0 ),
    .IQ(),
    .PAD(di[6])
  );

  defparam \di[5]_inst .imux.CONF = "1";
  defparam \di[5]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[5]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[5]_IN_to_TOP_I11_50_0 ),
    .IQ(),
    .PAD(di[5])
  );

  defparam \di[4]_inst .imux.CONF = "1";
  defparam \di[4]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[4]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[4]_IN_to_TOP_I21_53_0 ),
    .IQ(),
    .PAD(di[4])
  );

  defparam \di[3]_inst .imux.CONF = "1";
  defparam \di[3]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[3]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[3]_IN_to_TOP_I11_53_0 ),
    .IQ(),
    .PAD(di[3])
  );

  defparam \di[2]_inst .imux.CONF = "1";
  defparam \di[2]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[2]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[2]_IN_to_RIGHT_I14_54_0 ),
    .IQ(),
    .PAD(di[2])
  );

  defparam \di[1]_inst .imux.CONF = "1";
  defparam \di[1]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[1]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[1]_IN_to_RIGHT_I16_54_0 ),
    .IQ(),
    .PAD(di[1])
  );

  defparam \di[0]_inst .imux.CONF = "1";
  defparam \di[0]_inst .ioattrbox.CONF = "LVTTL";
  IOB \di[0]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-di[0]_IN_to_RIGHT_I18_54_0 ),
    .IQ(),
    .PAD(di[0])
  );

  defparam \do[15]_inst .driveattrbox.CONF = "12";
  defparam \do[15]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[15]_inst .omux.CONF = "O";
  defparam \do[15]_inst .outmux.CONF = "1";
  defparam \do[15]_inst .slew.CONF = "SLOW";
  IOB \do[15]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[15]_LEFT_O2_to_OUT17_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[15])
  );

  defparam \do[14]_inst .driveattrbox.CONF = "12";
  defparam \do[14]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[14]_inst .omux.CONF = "O";
  defparam \do[14]_inst .outmux.CONF = "1";
  defparam \do[14]_inst .slew.CONF = "SLOW";
  IOB \do[14]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[14]_LEFT_O2_to_OUT14_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[14])
  );

  defparam \do[13]_inst .driveattrbox.CONF = "12";
  defparam \do[13]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[13]_inst .omux.CONF = "O";
  defparam \do[13]_inst .outmux.CONF = "1";
  defparam \do[13]_inst .slew.CONF = "SLOW";
  IOB \do[13]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[13]_LEFT_O1_to_OUT16_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[13])
  );

  defparam \do[12]_inst .driveattrbox.CONF = "12";
  defparam \do[12]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[12]_inst .omux.CONF = "O";
  defparam \do[12]_inst .outmux.CONF = "1";
  defparam \do[12]_inst .slew.CONF = "SLOW";
  IOB \do[12]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[12]_LEFT_O2_to_OUT13_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[12])
  );

  defparam \do[11]_inst .driveattrbox.CONF = "12";
  defparam \do[11]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[11]_inst .omux.CONF = "O";
  defparam \do[11]_inst .outmux.CONF = "1";
  defparam \do[11]_inst .slew.CONF = "SLOW";
  IOB \do[11]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[11]_LEFT_O3_to_OUT13_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[11])
  );

  defparam \do[10]_inst .driveattrbox.CONF = "12";
  defparam \do[10]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[10]_inst .omux.CONF = "O";
  defparam \do[10]_inst .outmux.CONF = "1";
  defparam \do[10]_inst .slew.CONF = "SLOW";
  IOB \do[10]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[10]_LEFT_O1_to_OUT14_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[10])
  );

  defparam \do[9]_inst .driveattrbox.CONF = "12";
  defparam \do[9]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[9]_inst .omux.CONF = "O";
  defparam \do[9]_inst .outmux.CONF = "1";
  defparam \do[9]_inst .slew.CONF = "SLOW";
  IOB \do[9]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[9]_LEFT_O2_to_OUT9_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[9])
  );

  defparam \do[8]_inst .driveattrbox.CONF = "12";
  defparam \do[8]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[8]_inst .omux.CONF = "O";
  defparam \do[8]_inst .outmux.CONF = "1";
  defparam \do[8]_inst .slew.CONF = "SLOW";
  IOB \do[8]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[8]_LEFT_O3_to_OUT9_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[8])
  );

  defparam \do[7]_inst .driveattrbox.CONF = "12";
  defparam \do[7]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[7]_inst .omux.CONF = "O";
  defparam \do[7]_inst .outmux.CONF = "1";
  defparam \do[7]_inst .slew.CONF = "SLOW";
  IOB \do[7]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[7]_LEFT_O1_to_OUT10_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[7])
  );

  defparam \do[6]_inst .driveattrbox.CONF = "12";
  defparam \do[6]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[6]_inst .omux.CONF = "O";
  defparam \do[6]_inst .outmux.CONF = "1";
  defparam \do[6]_inst .slew.CONF = "SLOW";
  IOB \do[6]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[6]_LEFT_O2_to_OUT10_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[6])
  );

  defparam \do[5]_inst .driveattrbox.CONF = "12";
  defparam \do[5]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[5]_inst .omux.CONF = "O";
  defparam \do[5]_inst .outmux.CONF = "1";
  defparam \do[5]_inst .slew.CONF = "SLOW";
  IOB \do[5]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[5]_LEFT_O1_to_OUT8_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[5])
  );

  defparam \do[4]_inst .driveattrbox.CONF = "12";
  defparam \do[4]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[4]_inst .omux.CONF = "O";
  defparam \do[4]_inst .outmux.CONF = "1";
  defparam \do[4]_inst .slew.CONF = "SLOW";
  IOB \do[4]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[4]_LEFT_O1_to_OUT9_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[4])
  );

  defparam \do[3]_inst .driveattrbox.CONF = "12";
  defparam \do[3]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[3]_inst .omux.CONF = "O";
  defparam \do[3]_inst .outmux.CONF = "1";
  defparam \do[3]_inst .slew.CONF = "SLOW";
  IOB \do[3]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[3]_LEFT_O1_to_OUT4_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[3])
  );

  defparam \do[2]_inst .driveattrbox.CONF = "12";
  defparam \do[2]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[2]_inst .omux.CONF = "O";
  defparam \do[2]_inst .outmux.CONF = "1";
  defparam \do[2]_inst .slew.CONF = "SLOW";
  IOB \do[2]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[2]_LEFT_O3_to_OUT5_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[2])
  );

  defparam \do[1]_inst .driveattrbox.CONF = "12";
  defparam \do[1]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[1]_inst .omux.CONF = "O";
  defparam \do[1]_inst .outmux.CONF = "1";
  defparam \do[1]_inst .slew.CONF = "SLOW";
  IOB \do[1]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[1]_LEFT_O1_to_OUT6_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[1])
  );

  defparam \do[0]_inst .driveattrbox.CONF = "12";
  defparam \do[0]_inst .ioattrbox.CONF = "LVTTL";
  defparam \do[0]_inst .omux.CONF = "O";
  defparam \do[0]_inst .outmux.CONF = "1";
  defparam \do[0]_inst .slew.CONF = "SLOW";
  IOB \do[0]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_do_reg[0]_LEFT_O2_to_OUT6_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(do[0])
  );

  defparam rstn_inst.imux.CONF = "1";
  defparam rstn_inst.ioattrbox.CONF = "LVTTL";
  IOB rstn_inst (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-rstn_IN_to_RIGHT_I35_54_0 ),
    .IQ(),
    .PAD(rstn)
  );

  defparam iGclk_buf__0___inst.cemux.CONF = "1";
  defparam iGclk_buf__0___inst.disable_attr.CONF = "LOW";
  GCLK iGclk_buf__0___inst (
    .CE(),
    .IN(\net_Buf-pad-clk_CLKB_GCLKBUF1_IN_to_IN35_28_0 ),
    .OUT(\net_IBuf-clkpad-clk_OUT_to_CLKB_GCLK1_PW35_28_0 )
  );

  defparam clk_inst.ioattrbox.CONF = "LVTTL";
  GCLKIOB clk_inst (
    .PAD(clk),
    .GCLKOUT(\net_Buf-pad-clk_GCLKOUT_to_CLKB_CLKPAD135_28_0 )
  );

  defparam GSB_RHT_26_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_26_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_26_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_26_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_26_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_26_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_26_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_26_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llh11.CONF = "01";
  defparam GSB_RHT_26_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_26_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_26_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_26_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_26_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_26_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_26_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_26_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_26_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_26_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_26_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_26_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_26_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_26_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_26_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_26_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_26_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_26_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_26_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(\net_Buf-pad-di[15]_RIGHT_LLH11_to_LLH026_27_0 ),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(),
    .RIGHT_LLV6(),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(),
    .RIGHT_I3(\net_Buf-pad-di[15]_IN_to_RIGHT_I326_54_0 ),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_26_27_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_h6w1.CONF = "0001";
  defparam GSB_CNT_26_27_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_26_27_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_26_27_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_26_27_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_26_27_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_26_27_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_26_27_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_26_27_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_26_27_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_Buf-pad-di[15]_H6W1_to_H6E126_21_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_Buf-pad-di[15]_RIGHT_LLH11_to_LLH026_27_0 ),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_26_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_26_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_26_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_v6n2.CONF = "0101";
  defparam GSB_CNT_26_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_26_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_26_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_26_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_26_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_26_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_26_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(\net_Buf-pad-di[15]_H6W1_to_H6E126_21_0 ),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(\net_Buf-pad-di[15]_V6N2_to_V6S220_21_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_20_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_20_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_20_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_v6n2.CONF = "0000";
  defparam GSB_CNT_20_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_20_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_20_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_20_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_20_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_20_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_20_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(\net_Buf-pad-di[15]_V6N2_to_V6S213_21_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(\net_Buf-pad-di[15]_V6N2_to_V6S220_21_0 ),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_13_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_13_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_13_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_v6s1.CONF = "0101";
  defparam GSB_CNT_13_21_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n13.CONF = "01";
  defparam GSB_CNT_13_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n7.CONF = "01";
  defparam GSB_CNT_13_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_13_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_13_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_13_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_13_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_13_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_13_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(net_VCC_N7_to_S712_21_0),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(\net_Buf-pad-di[15]_N13_to_S1312_21_0 ),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(net_VCC_V6S1_to_V6N113_21_0),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(\net_Buf-pad-di[15]_V6N2_to_V6S213_21_0 ),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_12_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_llh0.CONF = "01";
  defparam GSB_CNT_12_21_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_12_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_12_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_12_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_out3.CONF = "001110";
  defparam GSB_CNT_12_21_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_out5.CONF = "001101";
  defparam GSB_CNT_12_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_12_21_0_inst.sps_s0_f_b1.CONF = "100110111";
  defparam GSB_CNT_12_21_0_inst.sps_s0_f_b2.CONF = "001111011";
  defparam GSB_CNT_12_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_21_0_inst.sps_s0_g_b1.CONF = "100101";
  defparam GSB_CNT_12_21_0_inst.sps_s0_g_b2.CONF = "001101";
  defparam GSB_CNT_12_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s0_sr_b.CONF = "110111";
  defparam GSB_CNT_12_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_12_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_12_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_12_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_12_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n12_e8.CONF = "0";
  defparam GSB_CNT_12_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_12_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_12_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(\net_Buf-pad-di[13]_W8_to_E812_21_0 ),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(\net_Buf-pad-di[13]_N12_to_S1211_21_0 ),
    .N13(),
    .N14(\net_Buf-pad-di[14]_S14_to_N1412_21_0 ),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(net_VCC_N7_to_S712_21_0),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(\net_Buf-pad-di[15]_N13_to_S1312_21_0 ),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[14]_LLH0_to_LLH012_8_0 ),
    .LLH6(\net_do_reg[15]_LLH6_to_LLH612_8_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK112_21_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(\net_Buf-pad-rstn_V6S1_to_V6D112_21_0 ),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-di[15]_S0_F_B1_to_F112_21_0 ),
    .S0_F_B2(net_VCC_S0_F_B2_to_F212_21_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Buf-pad-di[14]_S0_G_B1_to_G112_21_0 ),
    .S0_G_B2(net_VCC_S0_G_B2_to_G212_21_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK12_21_0 ),
    .S0_SR_B(\net_Buf-pad-rstn_S0_SR_B_to_SR12_21_0 ),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_do_reg[15]_XQ_to_S0_XQ12_21_0 ),
    .S0_YQ(\net_do_reg[14]_YQ_to_S0_YQ12_21_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_v6s1.CONF = "0000";
  defparam GSB_CNT_7_21_0_inst.sps_v6s2.CONF = "0000";
  defparam GSB_CNT_7_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n1.CONF = "10";
  defparam GSB_CNT_7_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n14.CONF = "0";
  defparam GSB_CNT_7_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_out0.CONF = "000111";
  defparam GSB_CNT_7_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_out2.CONF = "000111";
  defparam GSB_CNT_7_21_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_out4.CONF = "000111";
  defparam GSB_CNT_7_21_0_inst.sps_out5.CONF = "000111";
  defparam GSB_CNT_7_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_s13.CONF = "10";
  defparam GSB_CNT_7_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_s3.CONF = "01";
  defparam GSB_CNT_7_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s5.CONF = "01";
  defparam GSB_CNT_7_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_v6n7.CONF = "000";
  defparam GSB_CNT_7_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(net_VCC_N1_to_S16_21_0),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(net_VCC_N14_to_S146_21_0),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(\net_Buf-pad-di[8]_S3_to_N38_21_0 ),
    .S4(),
    .S5(\net_Buf-pad-di[9]_S5_to_N58_21_0 ),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(net_VCC_S13_to_N138_21_0),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(\net_Buf-pad-di[8]_H6W4_to_H6E47_21_0 ),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(net_VCC_V6N7_to_V6M74_21_0),
    .V6N8(\net_Buf-pad-di[9]_TOP_V6S8_to_V6N87_21_0 ),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(net_VCC_V6S1_to_V6N113_21_0),
    .V6S2(net_VCC_V6S2_to_V6M210_21_0),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(net_VCC_X_to_S0_X7_21_0),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_h6e2.CONF = "0010";
  defparam GSB_CNT_10_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s16.CONF = "01";
  defparam GSB_CNT_10_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_s22.CONF = "01";
  defparam GSB_CNT_10_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n18_e14.CONF = "0";
  defparam GSB_CNT_10_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(\net_Buf-pad-di[6]_W14_to_E1410_21_0 ),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(\net_Buf-pad-di[6]_N18_to_S189_21_0 ),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(net_VCC_S16_to_N1611_21_0),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(\net_Buf-pad-di[12]_S22_to_N2211_21_0 ),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(\net_Buf-pad-di[12]_V6S3_to_V6N310_21_0 ),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(net_VCC_V6S2_to_V6M210_21_0),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_llh0.CONF = "01";
  defparam GSB_CNT_11_21_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_11_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_v6s1.CONF = "0101";
  defparam GSB_CNT_11_21_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_out3.CONF = "001110";
  defparam GSB_CNT_11_21_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_out5.CONF = "001101";
  defparam GSB_CNT_11_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_11_21_0_inst.sps_s0_f_b1.CONF = "010111110";
  defparam GSB_CNT_11_21_0_inst.sps_s0_f_b2.CONF = "010101111";
  defparam GSB_CNT_11_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_21_0_inst.sps_s0_g_b1.CONF = "001010";
  defparam GSB_CNT_11_21_0_inst.sps_s0_g_b2.CONF = "010010";
  defparam GSB_CNT_11_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s0_sr_b.CONF = "001101";
  defparam GSB_CNT_11_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s14.CONF = "01";
  defparam GSB_CNT_11_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(net_VCC_S16_to_N1611_21_0),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(\net_Buf-pad-di[12]_S22_to_N2211_21_0 ),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(\net_Buf-pad-di[13]_N12_to_S1211_21_0 ),
    .S13(),
    .S14(\net_Buf-pad-di[14]_S14_to_N1412_21_0 ),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[12]_LLH0_to_LEFT_LLH611_2_0 ),
    .LLH6(\net_do_reg[13]_LLH6_to_LEFT_LLH011_2_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK111_21_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(\net_Buf-pad-rstn_V6S1_to_V6N111_21_0 ),
    .V6N2(\net_Buf-pad-di[14]_V6S2_to_V6N211_21_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(\net_Buf-pad-rstn_V6S1_to_V6D112_21_0 ),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-di[13]_S0_F_B1_to_F111_21_0 ),
    .S0_F_B2(net_VCC_S0_F_B2_to_F211_21_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Buf-pad-di[12]_S0_G_B1_to_G111_21_0 ),
    .S0_G_B2(net_VCC_S0_G_B2_to_G211_21_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK11_21_0 ),
    .S0_SR_B(\net_Buf-pad-rstn_S0_SR_B_to_SR11_21_0 ),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_do_reg[13]_XQ_to_S0_XQ11_21_0 ),
    .S0_YQ(\net_do_reg[12]_YQ_to_S0_YQ11_21_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_llh0.CONF = "01";
  defparam GSB_CNT_6_21_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_6_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_n9.CONF = "01";
  defparam GSB_CNT_6_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_out3.CONF = "001110";
  defparam GSB_CNT_6_21_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_out5.CONF = "001101";
  defparam GSB_CNT_6_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_6_21_0_inst.sps_s0_f_b1.CONF = "011011111";
  defparam GSB_CNT_6_21_0_inst.sps_s0_f_b2.CONF = "100111110";
  defparam GSB_CNT_6_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_21_0_inst.sps_s0_g_b1.CONF = "010100";
  defparam GSB_CNT_6_21_0_inst.sps_s0_g_b2.CONF = "100000";
  defparam GSB_CNT_6_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s0_sr_b.CONF = "110111";
  defparam GSB_CNT_6_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s17.CONF = "01";
  defparam GSB_CNT_6_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s5.CONF = "01";
  defparam GSB_CNT_6_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_v6s10.CONF = "101";
  defparam GSB_CNT_6_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s14_n14.CONF = "0";
  defparam GSB_CNT_6_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s17_n17.CONF = "0";
  defparam GSB_CNT_6_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s1_n1.CONF = "0";
  defparam GSB_CNT_6_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s5_n5.CONF = "0";
  defparam GSB_CNT_6_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(net_VCC_N1_to_S15_21_0),
    .N2(),
    .N3(),
    .N4(),
    .N5(\net_Buf-pad-di[4]_N5_to_S55_21_0 ),
    .N6(),
    .N7(),
    .N8(),
    .N9(\net_Buf-pad-di[11]_N9_to_S95_21_0 ),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(net_VCC_N14_to_S145_21_0),
    .N15(),
    .N16(),
    .N17(\net_Buf-pad-di[5]_N17_to_S175_21_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(\net_Buf-pad-di[0]_S23_to_N236_21_0 ),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(\net_Buf-pad-di[1]_E22_to_W226_21_0 ),
    .W23(),
    .S0(),
    .S1(net_VCC_N1_to_S16_21_0),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(net_VCC_N14_to_S146_21_0),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(\net_Buf-pad-di[11]_H6W8_to_H6E86_21_0 ),
    .H6E9(),
    .H6E10(\net_Buf-pad-di[7]_H6W10_to_H6E106_21_0 ),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[0]_LLH0_to_LEFT_LLH66_2_0 ),
    .LLH6(\net_do_reg[1]_LLH6_to_LEFT_LLH06_2_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK16_21_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(\net_Buf-pad-di[4]_TOP_V6D8_to_V6N86_21_0 ),
    .V6N9(),
    .V6N10(\net_Buf-pad-di[5]_TOP_V6D10_to_V6N106_21_0 ),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(\net_Buf-pad-di[7]_V6S10_to_V6M109_21_0 ),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(\net_Buf-pad-rstn_V6S1_to_V6N111_21_0 ),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-di[1]_S0_F_B1_to_F16_21_0 ),
    .S0_F_B2(net_VCC_S0_F_B2_to_F26_21_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Buf-pad-di[0]_S0_G_B1_to_G16_21_0 ),
    .S0_G_B2(net_VCC_S0_G_B2_to_G26_21_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK6_21_0 ),
    .S0_SR_B(\net_Buf-pad-rstn_S0_SR_B_to_SR6_21_0 ),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_do_reg[1]_XQ_to_S0_XQ6_21_0 ),
    .S0_YQ(\net_do_reg[0]_YQ_to_S0_YQ6_21_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_h6w2.CONF = "0010";
  defparam GSB_CNT_5_21_0_inst.sps_h6w3.CONF = "0001";
  defparam GSB_CNT_5_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_llh0.CONF = "00";
  defparam GSB_CNT_5_21_0_inst.sps_llh6.CONF = "00";
  defparam GSB_CNT_5_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_out7.CONF = "101011";
  defparam GSB_CNT_5_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_v6n1.CONF = "0100";
  defparam GSB_CNT_5_21_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_v6s1.CONF = "0011";
  defparam GSB_CNT_5_21_0_inst.sps_v6s2.CONF = "0101";
  defparam GSB_CNT_5_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_out2.CONF = "001101";
  defparam GSB_CNT_5_21_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_out4.CONF = "001110";
  defparam GSB_CNT_5_21_0_inst.sps_out5.CONF = "100111";
  defparam GSB_CNT_5_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_5_21_0_inst.sps_s0_f_b1.CONF = "001111101";
  defparam GSB_CNT_5_21_0_inst.sps_s0_f_b2.CONF = "100111110";
  defparam GSB_CNT_5_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_21_0_inst.sps_s0_g_b1.CONF = "100011";
  defparam GSB_CNT_5_21_0_inst.sps_s0_g_b2.CONF = "100000";
  defparam GSB_CNT_5_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_s0_sr_b.CONF = "001101";
  defparam GSB_CNT_5_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_s1_clk_b.CONF = "101011";
  defparam GSB_CNT_5_21_0_inst.sps_s1_f_b1.CONF = "011111110";
  defparam GSB_CNT_5_21_0_inst.sps_s1_f_b2.CONF = "010111011";
  defparam GSB_CNT_5_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_21_0_inst.sps_s1_g_b1.CONF = "100000";
  defparam GSB_CNT_5_21_0_inst.sps_s1_g_b2.CONF = "010101";
  defparam GSB_CNT_5_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_s1_sr_b.CONF = "001101";
  defparam GSB_CNT_5_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s23_w1.CONF = "0";
  defparam GSB_CNT_5_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(\net_Buf-pad-di[0]_E1_to_W15_21_0 ),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(\net_Buf-pad-di[10]_E9_to_W95_21_0 ),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(net_VCC_N1_to_S15_21_0),
    .S2(),
    .S3(),
    .S4(),
    .S5(\net_Buf-pad-di[4]_N5_to_S55_21_0 ),
    .S6(),
    .S7(),
    .S8(),
    .S9(\net_Buf-pad-di[11]_N9_to_S95_21_0 ),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(net_VCC_N14_to_S145_21_0),
    .S15(),
    .S16(),
    .S17(\net_Buf-pad-di[5]_N17_to_S175_21_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(\net_Buf-pad-di[0]_S23_to_N236_21_0 ),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(\net_Buf-pad-rstn_H6E1_to_H6M15_21_0 ),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(\net_do_reg[11]_H6W2_to_H6E25_14_0 ),
    .H6W3(\net_do_reg[10]_H6W3_to_H6E35_14_0 ),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[5]_LLH0_to_LLH05_8_0 ),
    .LLH6(\net_do_reg[4]_LLH6_to_LLH65_8_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK15_21_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(\net_Buf-pad-rstn_V6N1_to_V6A14_21_0 ),
    .V6N2(\net_Buf-pad-di[14]_TOP_V6C2_to_V6N25_21_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(\net_Buf-pad-rstn_V6S1_to_V6N111_21_0 ),
    .V6S2(\net_Buf-pad-di[14]_V6S2_to_V6N211_21_0 ),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-di[5]_S0_F_B1_to_F15_21_0 ),
    .S0_F_B2(net_VCC_S0_F_B2_to_F25_21_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Buf-pad-di[4]_S0_G_B1_to_G15_21_0 ),
    .S0_G_B2(net_VCC_S0_G_B2_to_G25_21_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK5_21_0 ),
    .S0_SR_B(\net_Buf-pad-rstn_S0_SR_B_to_SR5_21_0 ),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_do_reg[5]_XQ_to_S0_XQ5_21_0 ),
    .S0_YQ(\net_do_reg[4]_YQ_to_S0_YQ5_21_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Buf-pad-di[11]_S1_F_B1_to_F15_21_0 ),
    .S1_F_B2(net_VCC_S1_F_B2_to_F25_21_0),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(\net_Buf-pad-di[10]_S1_G_B1_to_G15_21_0 ),
    .S1_G_B2(net_VCC_S1_G_B2_to_G25_21_0),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK5_21_0 ),
    .S1_SR_B(\net_Buf-pad-rstn_S1_SR_B_to_SR5_21_0 ),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(\net_do_reg[11]_XQ_to_S1_XQ5_21_0 ),
    .S1_YQ(\net_do_reg[10]_YQ_to_S1_YQ5_21_0 ),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_llh0.CONF = "01";
  defparam GSB_CNT_8_21_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_8_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_out3.CONF = "101011";
  defparam GSB_CNT_8_21_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_out5.CONF = "100111";
  defparam GSB_CNT_8_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s1_clk_b.CONF = "101011";
  defparam GSB_CNT_8_21_0_inst.sps_s1_f_b1.CONF = "100111011";
  defparam GSB_CNT_8_21_0_inst.sps_s1_f_b2.CONF = "011111101";
  defparam GSB_CNT_8_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_21_0_inst.sps_s1_g_b1.CONF = "100100";
  defparam GSB_CNT_8_21_0_inst.sps_s1_g_b2.CONF = "011011";
  defparam GSB_CNT_8_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_s1_sr_b.CONF = "110111";
  defparam GSB_CNT_8_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s13_n13.CONF = "0";
  defparam GSB_CNT_8_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(\net_Buf-pad-di[8]_S3_to_N38_21_0 ),
    .N4(),
    .N5(\net_Buf-pad-di[9]_S5_to_N58_21_0 ),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(net_VCC_S13_to_N138_21_0),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(net_VCC_S13_to_N139_21_0),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[8]_LLH0_to_LLH08_8_0 ),
    .LLH6(\net_do_reg[9]_LLH6_to_LLH68_8_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK18_21_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_Buf-pad-rstn_V6S1_to_V6N111_21_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Buf-pad-di[9]_S1_F_B1_to_F18_21_0 ),
    .S1_F_B2(net_VCC_S1_F_B2_to_F28_21_0),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(\net_Buf-pad-di[8]_S1_G_B1_to_G18_21_0 ),
    .S1_G_B2(net_VCC_S1_G_B2_to_G28_21_0),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK8_21_0 ),
    .S1_SR_B(\net_Buf-pad-rstn_S1_SR_B_to_SR8_21_0 ),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(\net_do_reg[9]_XQ_to_S1_XQ8_21_0 ),
    .S1_YQ(\net_do_reg[8]_YQ_to_S1_YQ8_21_0 ),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_llh0.CONF = "01";
  defparam GSB_CNT_9_21_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_9_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_w1.CONF = "0";
  defparam GSB_CNT_9_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_out3.CONF = "101011";
  defparam GSB_CNT_9_21_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_out5.CONF = "100111";
  defparam GSB_CNT_9_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s1_clk_b.CONF = "101011";
  defparam GSB_CNT_9_21_0_inst.sps_s1_f_b1.CONF = "100101111";
  defparam GSB_CNT_9_21_0_inst.sps_s1_f_b2.CONF = "011111101";
  defparam GSB_CNT_9_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_21_0_inst.sps_s1_g_b1.CONF = "011011";
  defparam GSB_CNT_9_21_0_inst.sps_s1_g_b2.CONF = "011011";
  defparam GSB_CNT_9_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_s1_sr_b.CONF = "111011";
  defparam GSB_CNT_9_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(net_VCC_S13_to_N139_21_0),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(\net_Buf-pad-di[6]_N18_to_S189_21_0 ),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[6]_LLH0_to_LEFT_LLH69_2_0 ),
    .LLH6(\net_do_reg[7]_LLH6_to_LEFT_LLH09_2_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK19_21_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(\net_Buf-pad-di[7]_V6S10_to_V6M109_21_0 ),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(\net_Buf-pad-rstn_V6S1_to_V6N111_21_0 ),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Buf-pad-di[7]_S1_F_B1_to_F19_21_0 ),
    .S1_F_B2(net_VCC_S1_F_B2_to_F29_21_0),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(\net_Buf-pad-di[6]_S1_G_B1_to_G19_21_0 ),
    .S1_G_B2(net_VCC_S1_G_B2_to_G29_21_0),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK9_21_0 ),
    .S1_SR_B(\net_Buf-pad-rstn_S1_SR_B_to_SR9_21_0 ),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(\net_do_reg[7]_XQ_to_S1_XQ9_21_0 ),
    .S1_YQ(\net_do_reg[6]_YQ_to_S1_YQ9_21_0 ),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_21_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_llh0.CONF = "01";
  defparam GSB_CNT_4_21_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_4_21_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_21_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_21_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_v6s3.CONF = "0100";
  defparam GSB_CNT_4_21_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w12.CONF = "0";
  defparam GSB_CNT_4_21_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e12.CONF = "10";
  defparam GSB_CNT_4_21_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_out3.CONF = "001101";
  defparam GSB_CNT_4_21_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_out5.CONF = "001110";
  defparam GSB_CNT_4_21_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_4_21_0_inst.sps_s0_f_b1.CONF = "010110111";
  defparam GSB_CNT_4_21_0_inst.sps_s0_f_b2.CONF = "001110111";
  defparam GSB_CNT_4_21_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_21_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_21_0_inst.sps_s0_g_b1.CONF = "011100";
  defparam GSB_CNT_4_21_0_inst.sps_s0_g_b2.CONF = "001111";
  defparam GSB_CNT_4_21_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s0_sr_b.CONF = "101101";
  defparam GSB_CNT_4_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_21_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_21_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_21_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_21_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_21_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_21_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(\net_Buf-pad-di[2]_E22_to_W224_21_0 ),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(\net_Buf-pad-di[12]_H6W2_to_H6E24_21_0 ),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[3]_LLH0_to_LLH04_8_0 ),
    .LLH6(\net_do_reg[2]_LLH6_to_LEFT_LLH04_2_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK14_21_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(\net_Buf-pad-di[3]_TOP_V6S6_to_V6M64_21_0 ),
    .V6M7(net_VCC_V6N7_to_V6M74_21_0),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(\net_Buf-pad-di[12]_V6S3_to_V6N310_21_0 ),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(\net_Buf-pad-rstn_V6N1_to_V6A14_21_0 ),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-di[3]_S0_F_B1_to_F14_21_0 ),
    .S0_F_B2(net_VCC_S0_F_B2_to_F24_21_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Buf-pad-di[2]_S0_G_B1_to_G14_21_0 ),
    .S0_G_B2(net_VCC_S0_G_B2_to_G24_21_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK4_21_0 ),
    .S0_SR_B(\net_Buf-pad-rstn_S0_SR_B_to_SR4_21_0 ),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_do_reg[3]_XQ_to_S0_XQ4_21_0 ),
    .S0_YQ(\net_do_reg[2]_YQ_to_S0_YQ4_21_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_21_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w2.CONF = "00111011";
  defparam GSB_TOP_1_21_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_21_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_21_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6e1.CONF = "00111011";
  defparam GSB_TOP_1_21_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s6.CONF = "111011";
  defparam GSB_TOP_1_21_0_inst.sps_v6s8.CONF = "110111";
  defparam GSB_TOP_1_21_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6c2.CONF = "01110";
  defparam GSB_TOP_1_21_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d10.CONF = "110111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d8.CONF = "111011";
  defparam GSB_TOP_1_21_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_21_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(\net_Buf-pad-di[5]_TOP_H6E2_to_TOP_H6M21_21_0 ),
    .TOP_H6M3(\net_Buf-pad-di[9]_TOP_H6W3_to_TOP_H6M31_21_0 ),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(\net_Buf-pad-di[14]_TOP_V6C2_to_V6N25_21_0 ),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(\net_Buf-pad-di[4]_TOP_V6D8_to_V6N86_21_0 ),
    .TOP_V6D9(),
    .TOP_V6D10(\net_Buf-pad-di[5]_TOP_V6D10_to_V6N106_21_0 ),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(\net_Buf-pad-di[3]_TOP_V6S6_to_V6M64_21_0 ),
    .TOP_V6S7(),
    .TOP_V6S8(\net_Buf-pad-di[9]_TOP_V6S8_to_V6N87_21_0 ),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(\net_Buf-pad-di[3]_TOP_LLH6_to_TOP_LLH01_21_0 ),
    .TOP_LLH6(\net_Buf-pad-di[4]_TOP_LLH0_to_TOP_LLH61_21_0 ),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(\net_Buf-pad-di[14]_IN_to_TOP_I11_21_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_35_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w0.CONF = "01011011";
  defparam GSB_TOP_1_35_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_35_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_35_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_35_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(\net_Buf-pad-di[13]_TOP_H6W0_to_TOP_H6E01_29_0 ),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(\net_Buf-pad-di[13]_IN_to_TOP_I11_35_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_29_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6w0.CONF = "01101110";
  defparam GSB_TOP_1_29_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_29_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_29_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_29_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_29_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_29_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_29_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_29_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(\net_Buf-pad-di[13]_TOP_H6W0_to_TOP_H6E01_29_0 ),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(\net_Buf-pad-di[13]_TOP_H6W0_to_TOP_H6E01_22_0 ),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_22_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6w3.CONF = "00111011";
  defparam GSB_TOP_1_22_0_inst.sps_h6w4.CONF = "01101110";
  defparam GSB_TOP_1_22_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_22_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_22_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_22_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_22_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_22_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_v6s6.CONF = "101111";
  defparam GSB_TOP_1_22_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_22_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_22_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_22_0_inst.sps_v6d8.CONF = "101111";
  defparam GSB_TOP_1_22_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_22_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_22_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(\net_Buf-pad-di[13]_TOP_H6W0_to_TOP_H6E01_22_0 ),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(\net_Buf-pad-di[10]_TOP_H6W4_to_TOP_H6C41_20_0 ),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(\net_Buf-pad-di[13]_TOP_V6D8_to_V6N86_22_0 ),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(\net_Buf-pad-di[6]_TOP_V6S6_to_V6N67_22_0 ),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(\net_Buf-pad-di[10]_TOP_LLH6_to_TOP_LLH01_22_0 ),
    .TOP_LLH6(\net_Buf-pad-di[6]_TOP_LLH6_to_TOP_LLH61_22_0 ),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_CNT_6_22_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_22_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_22_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_22_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_22_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_22_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_22_0_inst.sps_v6s8.CONF = "000";
  defparam GSB_CNT_6_22_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_22_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_22_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(\net_Buf-pad-di[13]_TOP_V6D8_to_V6N86_22_0 ),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(\net_Buf-pad-di[13]_V6S8_to_V6N812_22_0 ),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_12_22_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_12_22_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_12_22_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_w8.CONF = "10";
  defparam GSB_CNT_12_22_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_12_22_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_12_22_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_12_22_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_12_22_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_12_22_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_12_22_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(\net_Buf-pad-di[13]_W8_to_E812_21_0 ),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(\net_Buf-pad-di[13]_V6S8_to_V6N812_22_0 ),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_40_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6w1.CONF = "01101110";
  defparam GSB_TOP_1_40_0_inst.sps_h6w2.CONF = "01011011";
  defparam GSB_TOP_1_40_0_inst.sps_h6w3.CONF = "01011110";
  defparam GSB_TOP_1_40_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_40_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_40_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_v6s10.CONF = "101111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_40_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(\net_Buf-pad-di[7]_TOP_H6W1_to_TOP_H6E11_40_0 ),
    .TOP_H6E2(),
    .TOP_H6E3(\net_Buf-pad-di[8]_TOP_H6W3_to_TOP_H6E31_40_0 ),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(\net_Buf-pad-di[7]_TOP_H6W1_to_TOP_H6E11_34_0 ),
    .TOP_H6W2(\net_Buf-pad-di[11]_TOP_H6W2_to_TOP_H6E21_34_0 ),
    .TOP_H6W3(\net_Buf-pad-di[12]_TOP_H6W3_to_TOP_H6E31_34_0 ),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(\net_Buf-pad-di[8]_TOP_V6S10_to_V6N107_40_0 ),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(\net_Buf-pad-di[12]_IN_to_TOP_I21_40_0 ),
    .TOP_I1(\net_Buf-pad-di[11]_IN_to_TOP_I11_40_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_34_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6w1.CONF = "01101110";
  defparam GSB_TOP_1_34_0_inst.sps_h6w2.CONF = "01101110";
  defparam GSB_TOP_1_34_0_inst.sps_h6w3.CONF = "01101110";
  defparam GSB_TOP_1_34_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_34_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_34_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_34_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(\net_Buf-pad-di[7]_TOP_H6W1_to_TOP_H6E11_34_0 ),
    .TOP_H6E2(\net_Buf-pad-di[11]_TOP_H6W2_to_TOP_H6E21_34_0 ),
    .TOP_H6E3(\net_Buf-pad-di[12]_TOP_H6W3_to_TOP_H6E31_34_0 ),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(\net_Buf-pad-di[7]_TOP_H6W1_to_TOP_H6E11_27_0 ),
    .TOP_H6W2(\net_Buf-pad-di[11]_TOP_H6W2_to_TOP_H6E21_27_0 ),
    .TOP_H6W3(\net_Buf-pad-di[12]_TOP_H6W3_to_TOP_H6E31_27_0 ),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_27_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_27_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_27_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s2.CONF = "0011111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d4.CONF = "101111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d6.CONF = "111011";
  defparam GSB_TOP_1_27_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_27_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(\net_Buf-pad-di[7]_TOP_H6W1_to_TOP_H6E11_27_0 ),
    .TOP_H6E2(\net_Buf-pad-di[11]_TOP_H6W2_to_TOP_H6E21_27_0 ),
    .TOP_H6E3(\net_Buf-pad-di[12]_TOP_H6W3_to_TOP_H6E31_27_0 ),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(\net_Buf-pad-di[11]_TOP_V6D4_to_V6N46_27_0 ),
    .TOP_V6D5(),
    .TOP_V6D6(\net_Buf-pad-di[7]_TOP_V6D6_to_V6N66_27_0 ),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(\net_Buf-pad-di[12]_TOP_V6S2_to_V6M24_27_0 ),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_CNT_4_27_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_h6w2.CONF = "0011";
  defparam GSB_CNT_4_27_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_27_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_27_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_27_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_27_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_27_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_27_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_27_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_27_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(\net_Buf-pad-di[12]_H6W2_to_H6E24_21_0 ),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(\net_Buf-pad-di[12]_TOP_V6S2_to_V6M24_27_0 ),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_27_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_h6w10.CONF = "011";
  defparam GSB_CNT_6_27_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_h6w8.CONF = "011";
  defparam GSB_CNT_6_27_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_27_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_27_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_27_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_27_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_27_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_27_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_27_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_27_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(\net_Buf-pad-di[11]_H6W8_to_H6E86_21_0 ),
    .H6W9(),
    .H6W10(\net_Buf-pad-di[7]_H6W10_to_H6E106_21_0 ),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(\net_Buf-pad-di[11]_TOP_V6D4_to_V6N46_27_0 ),
    .V6N5(),
    .V6N6(\net_Buf-pad-di[7]_TOP_V6D6_to_V6N66_27_0 ),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_42_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_42_0_inst.sps_llh6.CONF = "0111011111";
  defparam GSB_TOP_1_42_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_42_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(\net_Buf-pad-di[10]_TOP_LLH6_to_TOP_LLH01_22_0 ),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(\net_Buf-pad-di[10]_IN_to_TOP_I21_42_0 ),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_20_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_20_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_20_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_20_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_llv8.CONF = "00";
  defparam GSB_TOP_1_20_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_20_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_20_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_20_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_20_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(\net_Buf-pad-di[10]_TOP_H6W4_to_TOP_H6C41_20_0 ),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(\net_Buf-pad-di[10]_TOP_LLV8_to_LLV05_20_0 ),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_CNT_5_20_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_20_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_20_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_v6n1.CONF = "0010";
  defparam GSB_CNT_5_20_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e1.CONF = "01";
  defparam GSB_CNT_5_20_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_e9.CONF = "10";
  defparam GSB_CNT_5_20_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_20_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_20_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_20_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_20_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_20_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_20_0_inst (
    .E0(),
    .E1(\net_Buf-pad-di[0]_E1_to_W15_21_0 ),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(\net_Buf-pad-di[10]_E9_to_W95_21_0 ),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(\net_Buf-pad-di[0]_V6N0_to_V6M05_20_0 ),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(\net_Buf-pad-di[10]_TOP_LLV8_to_LLV05_20_0 ),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_44_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_llh0.CONF = "0111110111";
  defparam GSB_TOP_1_44_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_44_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_44_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(\net_Buf-pad-di[9]_TOP_LLH0_to_TOP_LLH61_24_0 ),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(\net_Buf-pad-di[9]_IN_to_TOP_I11_44_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_24_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6w3.CONF = "00111011";
  defparam GSB_TOP_1_24_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_24_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_24_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_24_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_24_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_24_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_24_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_24_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(\net_Buf-pad-di[9]_TOP_H6W3_to_TOP_H6M31_21_0 ),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(\net_Buf-pad-di[9]_TOP_LLH0_to_TOP_LLH61_24_0 ),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_47_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6w1.CONF = "01011011";
  defparam GSB_TOP_1_47_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6w3.CONF = "01011110";
  defparam GSB_TOP_1_47_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_47_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_47_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_47_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(\net_Buf-pad-di[7]_TOP_H6W1_to_TOP_H6E11_40_0 ),
    .TOP_H6W2(),
    .TOP_H6W3(\net_Buf-pad-di[8]_TOP_H6W3_to_TOP_H6E31_40_0 ),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(\net_Buf-pad-di[8]_IN_to_TOP_I21_47_0 ),
    .TOP_I1(\net_Buf-pad-di[7]_IN_to_TOP_I11_47_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_CNT_7_40_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_h6w4.CONF = "011";
  defparam GSB_CNT_7_40_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_40_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_40_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_40_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_40_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_40_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_40_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_40_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_40_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(\net_Buf-pad-di[8]_H6W4_to_H6E47_34_0 ),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(\net_Buf-pad-di[8]_TOP_V6S10_to_V6N107_40_0 ),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_34_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_h6w4.CONF = "101";
  defparam GSB_CNT_7_34_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_34_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_34_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_34_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_34_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_34_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_34_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_34_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_34_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(\net_Buf-pad-di[8]_H6W4_to_H6E47_34_0 ),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(\net_Buf-pad-di[8]_H6W4_to_H6E47_27_0 ),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_27_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_h6w4.CONF = "101";
  defparam GSB_CNT_7_27_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_27_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_27_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_27_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_27_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_27_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_27_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_27_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_27_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(\net_Buf-pad-di[8]_H6W4_to_H6E47_27_0 ),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(\net_Buf-pad-di[8]_H6W4_to_H6E47_21_0 ),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_48_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_48_0_inst.sps_llh6.CONF = "0111011111";
  defparam GSB_TOP_1_48_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_48_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(\net_Buf-pad-di[6]_TOP_LLH6_to_TOP_LLH61_22_0 ),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(\net_Buf-pad-di[6]_IN_to_TOP_I21_48_0 ),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_CNT_7_22_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_22_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_22_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_22_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_22_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_22_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.sps_v6s6.CONF = "000";
  defparam GSB_CNT_7_22_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_22_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_22_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_22_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(\net_Buf-pad-di[6]_TOP_V6S6_to_V6N67_22_0 ),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(\net_Buf-pad-di[6]_V6S6_to_V6M610_22_0 ),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_22_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_22_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_22_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_w14.CONF = "0";
  defparam GSB_CNT_10_22_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_22_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_22_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_22_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_22_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_22_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_22_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(\net_Buf-pad-di[6]_W14_to_E1410_21_0 ),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(\net_Buf-pad-di[6]_V6S6_to_V6M610_22_0 ),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_50_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_llh0.CONF = "0111110111";
  defparam GSB_TOP_1_50_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_50_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_50_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(\net_Buf-pad-di[5]_TOP_LLH0_to_TOP_LLH61_18_0 ),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(\net_Buf-pad-di[5]_IN_to_TOP_I11_50_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_18_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_18_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_18_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6e2.CONF = "00111011";
  defparam GSB_TOP_1_18_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_18_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_18_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_18_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_18_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_18_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(\net_Buf-pad-di[5]_TOP_H6E2_to_TOP_H6M21_21_0 ),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(\net_Buf-pad-di[5]_TOP_LLH0_to_TOP_LLH61_18_0 ),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_53_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_llh0.CONF = "0111011111";
  defparam GSB_TOP_1_53_0_inst.sps_llh6.CONF = "0111110111";
  defparam GSB_TOP_1_53_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_53_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(\net_Buf-pad-di[4]_TOP_LLH0_to_TOP_LLH61_21_0 ),
    .TOP_LLH6(\net_Buf-pad-di[3]_TOP_LLH6_to_TOP_LLH01_21_0 ),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(\net_Buf-pad-di[4]_IN_to_TOP_I21_53_0 ),
    .TOP_I1(\net_Buf-pad-di[3]_IN_to_TOP_I11_53_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_RHT_4_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_4_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_4_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_4_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_4_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh4.CONF = "00";
  defparam GSB_RHT_4_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_4_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_4_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_4_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_4_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_4_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_4_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_4_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_4_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(\net_Buf-pad-di[2]_RIGHT_LLH4_to_LLH04_20_0 ),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(),
    .RIGHT_LLV6(),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(\net_Buf-pad-di[2]_IN_to_RIGHT_I14_54_0 ),
    .RIGHT_I2(),
    .RIGHT_I3(),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_4_20_0_inst.sps_h6w0.CONF = "0001";
  defparam GSB_CNT_4_20_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_20_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_20_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e22.CONF = "10";
  defparam GSB_CNT_4_20_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_20_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_20_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_20_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_20_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_20_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_20_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(\net_Buf-pad-di[2]_E22_to_W224_21_0 ),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_Buf-pad-di[2]_RIGHT_LLH4_to_LLH04_20_0 ),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_RHT_6_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_6_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_6_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_6_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_6_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh4.CONF = "00";
  defparam GSB_RHT_6_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_6_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_6_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_6_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_6_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_6_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_6_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_6_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_6_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(\net_Buf-pad-di[1]_RIGHT_LLH4_to_LLH06_20_0 ),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(),
    .RIGHT_LLV6(),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(\net_Buf-pad-di[1]_IN_to_RIGHT_I16_54_0 ),
    .RIGHT_I2(),
    .RIGHT_I3(),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_6_20_0_inst.sps_h6w0.CONF = "0001";
  defparam GSB_CNT_6_20_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_20_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_20_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e22.CONF = "10";
  defparam GSB_CNT_6_20_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_20_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_20_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_20_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_20_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_20_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_20_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(\net_Buf-pad-di[1]_E22_to_W226_21_0 ),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_Buf-pad-di[1]_RIGHT_LLH4_to_LLH06_20_0 ),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_RHT_8_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_8_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_8_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_8_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_8_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh4.CONF = "00";
  defparam GSB_RHT_8_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_8_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_8_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_8_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_8_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_8_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_8_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_8_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_8_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(\net_Buf-pad-di[0]_RIGHT_LLH4_to_LLH08_20_0 ),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(),
    .RIGHT_LLV6(),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(\net_Buf-pad-di[0]_IN_to_RIGHT_I18_54_0 ),
    .RIGHT_I2(),
    .RIGHT_I3(),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_8_20_0_inst.sps_h6w0.CONF = "0001";
  defparam GSB_CNT_8_20_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_20_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_20_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_v6n0.CONF = "0011";
  defparam GSB_CNT_8_20_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_20_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_20_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_20_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_20_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_20_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_20_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_Buf-pad-di[0]_RIGHT_LLH4_to_LLH08_20_0 ),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(\net_Buf-pad-di[0]_V6N0_to_V6M05_20_0 ),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CLKB_35_28_0_inst.sps_h6d0.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6d1.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6d2.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6d3.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh1.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh10.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh4.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh7.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e0.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e1.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e2.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e3.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.spbu_gclk0.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_gclk1.CONF = "0";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e0.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e1.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e2.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e3.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w0.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w1.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w2.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w3.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.sps_ce0.CONF = "1111";
  defparam GSB_CLKB_35_28_0_inst.sps_ce1.CONF = "1111";
  defparam GSB_CLKB_35_28_0_inst.sps_clkfbl.CONF = "010";
  defparam GSB_CLKB_35_28_0_inst.sps_clkfbr.CONF = "010";
  defparam GSB_CLKB_35_28_0_inst.sps_clkinl.CONF = "011";
  defparam GSB_CLKB_35_28_0_inst.sps_clkinr.CONF = "011";
  defparam GSB_CLKB_35_28_0_inst.sps_gclkbuf0_in.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_gclkbuf1_in.CONF = "011111";
  GSB_CLKB GSB_CLKB_35_28_0_inst (
    .CLKB_H6E0(),
    .CLKB_H6E1(),
    .CLKB_H6E2(),
    .CLKB_H6E3(),
    .CLKB_H6A0(),
    .CLKB_H6A1(),
    .CLKB_H6A2(),
    .CLKB_H6A3(),
    .CLKB_H6B0(),
    .CLKB_H6B1(),
    .CLKB_H6B2(),
    .CLKB_H6B3(),
    .CLKB_H6M0(),
    .CLKB_H6M1(),
    .CLKB_H6M2(),
    .CLKB_H6M3(),
    .CLKB_H6C0(),
    .CLKB_H6C1(),
    .CLKB_H6C2(),
    .CLKB_H6C3(),
    .CLKB_H6D0(),
    .CLKB_H6D1(),
    .CLKB_H6D2(),
    .CLKB_H6D3(),
    .CLKB_LLH1(),
    .CLKB_LLH4(),
    .CLKB_LLH7(),
    .CLKB_LLH10(),
    .CLKB_GCLK0(),
    .CLKB_GCLK1(\net_IBuf-clkpad-clk_CLKB_GCLK1_to_CLKC_GCLK118_28_0 ),
    .CLKB_VGCLK0(),
    .CLKB_VGCLK1(),
    .CLKB_VGCLK2(),
    .CLKB_VGCLK3(),
    .CLKB_HGCLK_E0(),
    .CLKB_HGCLK_E1(),
    .CLKB_HGCLK_E2(),
    .CLKB_HGCLK_E3(),
    .CLKB_HGCLK_W0(),
    .CLKB_HGCLK_W1(),
    .CLKB_HGCLK_W2(),
    .CLKB_HGCLK_W3(),
    .CLKB_CLKINL_1(),
    .CLKB_CLKFBL_1(),
    .CLKB_CLKDVL_1(),
    .CLKB_CLK0L_1(),
    .CLKB_CLK90L_1(),
    .CLKB_CLK180L_1(),
    .CLKB_CLK270L_1(),
    .CLKB_CLK2XL_1(),
    .CLKB_CLK2X90L_1(),
    .CLKB_LOCKEDL_1(),
    .CLKB_CLKINR_1(),
    .CLKB_CLKFBR_1(),
    .CLKB_CLKDVR_1(),
    .CLKB_CLK0R_1(),
    .CLKB_CLK90R_1(),
    .CLKB_CLK180R_1(),
    .CLKB_CLK270R_1(),
    .CLKB_CLK2XR_1(),
    .CLKB_CLK2X90R_1(),
    .CLKB_LOCKEDR_1(),
    .CLKB_CLKPAD0(),
    .CLKB_CLKPAD1(\net_Buf-pad-clk_GCLKOUT_to_CLKB_CLKPAD135_28_0 ),
    .CLKB_GCLKBUF0_IN(),
    .CLKB_GCLK0_PW(),
    .CLKB_CE0(),
    .CLKB_GCLKBUF1_IN(\net_Buf-pad-clk_CLKB_GCLKBUF1_IN_to_IN35_28_0 ),
    .CLKB_GCLK1_PW(\net_IBuf-clkpad-clk_OUT_to_CLKB_GCLK1_PW35_28_0 ),
    .CLKB_CE1(),
    .BOT_CLKINL(),
    .BOT_CLKFBL(),
    .BOT_CLKINR(),
    .BOT_CLKFBR(),
    .DLL1_RST_I(),
    .DLL1_RST_O(),
    .DLL0_RST_I(),
    .DLL0_RST_O()
  );

  defparam GSB_CNT_12_8_0_inst.sps_h6w0.CONF = "0001";
  defparam GSB_CNT_12_8_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w3.CONF = "0000";
  defparam GSB_CNT_12_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_12_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_12_8_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_12_8_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(\net_do_reg[14]_H6W0_to_LEFT_H6E012_2_0 ),
    .H6W1(),
    .H6W2(),
    .H6W3(\net_do_reg[15]_H6W3_to_LEFT_H6E312_2_0 ),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[14]_LLH0_to_LLH012_8_0 ),
    .LLH6(\net_do_reg[15]_LLH6_to_LLH612_8_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_12_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_12_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_12_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_12_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_12_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_12_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_12_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_12_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_12_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_12_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_12_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_12_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_12_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_12_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_12_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_12_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_12_2_0_inst.sps_v6s0.CONF = "00111110";
  defparam GSB_LFT_12_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_12_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_12_2_0_inst.sps_v6s3.CONF = "00111110";
  defparam GSB_LFT_12_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_12_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_12_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_12_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_12_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_12_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_12_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_12_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_12_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_12_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_12_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_12_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_12_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_12_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_12_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_12_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(\net_do_reg[14]_H6W0_to_LEFT_H6E012_2_0 ),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(\net_do_reg[15]_H6W3_to_LEFT_H6E312_2_0 ),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(\net_do_reg[14]_LEFT_V6S0_to_LEFT_V6M015_2_0 ),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(\net_do_reg[15]_LEFT_V6S3_to_LEFT_V6N319_2_0 ),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_LFT_19_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_19_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_19_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_19_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_19_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_19_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_19_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_19_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_19_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_19_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_19_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_19_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_19_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_19_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_19_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_19_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e20.CONF = "01";
  defparam GSB_LFT_19_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_19_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_19_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_19_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_19_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_19_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_19_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_19_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_19_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_19_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_19_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_19_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(\net_do_reg[15]_LEFT_E20_to_W2019_3_0 ),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(\net_do_reg[15]_LEFT_V6S3_to_LEFT_V6N319_2_0 ),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_19_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_19_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_19_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_19_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_19_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_19_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_19_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n19_w20.CONF = "0";
  defparam GSB_CNT_19_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_19_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_19_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(\net_do_reg[15]_N19_to_S1917_3_0 ),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(\net_do_reg[15]_LEFT_E20_to_W2019_3_0 ),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_17_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_17_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_17_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_17_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_17_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_17_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_17_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n1_w2.CONF = "0";
  defparam GSB_CNT_17_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s19_w21.CONF = "0";
  defparam GSB_CNT_17_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_17_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_17_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(\net_do_reg[13]_N1_to_S116_3_0 ),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(\net_do_reg[13]_LEFT_E2_to_W217_3_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(\net_do_reg[15]_W21_to_LEFT_E2117_2_0 ),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(\net_do_reg[15]_N19_to_S1917_3_0 ),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_17_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_17_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_17_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_17_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_17_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_17_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_17_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_17_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_17_2_0_inst.sps_o2.CONF = "110001011";
  defparam GSB_LFT_17_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_17_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_17_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_17_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_17_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_17_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_17_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e2.CONF = "01";
  defparam GSB_LFT_17_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_17_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_17_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_17_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_17_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_17_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_17_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_17_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_17_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_17_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_17_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_17_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(\net_do_reg[15]_W21_to_LEFT_E2117_2_0 ),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(\net_do_reg[13]_LEFT_E2_to_W217_3_0 ),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(\net_do_reg[13]_LEFT_V6S0_to_LEFT_V6N017_2_0 ),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(\net_do_reg[15]_LEFT_O2_to_OUT17_2_0 ),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_LFT_15_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_15_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_15_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_15_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_15_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_15_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_15_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_15_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_15_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_15_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_15_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_15_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_15_2_0_inst.sps_e1.CONF = "01";
  defparam GSB_LFT_15_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_15_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_15_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_15_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_15_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_15_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_15_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_15_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_15_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_15_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_15_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_15_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_15_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_15_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_15_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(\net_do_reg[14]_LEFT_E1_to_W115_3_0 ),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(\net_do_reg[14]_LEFT_V6S0_to_LEFT_V6M015_2_0 ),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_15_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_15_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_15_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_15_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_15_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_15_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_15_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n20_w1.CONF = "0";
  defparam GSB_CNT_15_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_15_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_15_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(\net_do_reg[14]_N20_to_S2014_3_0 ),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(\net_do_reg[14]_LEFT_E1_to_W115_3_0 ),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_14_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_14_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_14_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n14_w19.CONF = "0";
  defparam GSB_CNT_14_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n15_w16.CONF = "0";
  defparam GSB_CNT_14_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s20_w22.CONF = "0";
  defparam GSB_CNT_14_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_14_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(\net_do_reg[12]_N14_to_S1413_3_0 ),
    .N15(\net_do_reg[11]_N15_to_S1513_3_0 ),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(\net_do_reg[11]_LEFT_E16_to_W1614_3_0 ),
    .W17(),
    .W18(),
    .W19(\net_do_reg[12]_LEFT_E19_to_W1914_3_0 ),
    .W20(),
    .W21(),
    .W22(\net_do_reg[14]_W22_to_LEFT_E2214_2_0 ),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(\net_do_reg[14]_N20_to_S2014_3_0 ),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_14_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_14_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_14_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_14_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_14_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_14_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_14_2_0_inst.sps_o1.CONF = "110111110";
  defparam GSB_LFT_14_2_0_inst.sps_o2.CONF = "110001101";
  defparam GSB_LFT_14_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_14_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e16.CONF = "01";
  defparam GSB_LFT_14_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e19.CONF = "01";
  defparam GSB_LFT_14_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_14_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_14_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(\net_do_reg[14]_W22_to_LEFT_E2214_2_0 ),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(\net_do_reg[12]_LEFT_E19_to_W1914_3_0 ),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(\net_do_reg[11]_LEFT_E16_to_W1614_3_0 ),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(\net_do_reg[10]_H6W1_to_LEFT_H6E114_2_0 ),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(\net_do_reg[11]_LEFT_V6S2_to_LEFT_V6M214_2_0 ),
    .LEFT_V6M3(\net_do_reg[12]_LEFT_V6S3_to_LEFT_V6M314_2_0 ),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_do_reg[10]_LEFT_O1_to_OUT14_2_0 ),
    .LEFT_O2(\net_do_reg[14]_LEFT_O2_to_OUT14_2_0 ),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_LFT_11_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_11_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_11_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_11_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_11_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_11_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_11_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_11_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_11_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_11_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6s0.CONF = "00111110";
  defparam GSB_LFT_11_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6s2.CONF = "01101110";
  defparam GSB_LFT_11_2_0_inst.sps_v6s3.CONF = "00111110";
  defparam GSB_LFT_11_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e0.CONF = "0111011";
  defparam GSB_LFT_11_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e3.CONF = "0111011";
  defparam GSB_LFT_11_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_11_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_11_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(\net_do_reg[13]_LLH6_to_LEFT_LLH011_2_0 ),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(\net_do_reg[12]_LLH0_to_LEFT_LLH611_2_0 ),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(\net_do_reg[11]_LEFT_V6S2_to_LEFT_V6N211_2_0 ),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(\net_do_reg[13]_LEFT_V6S0_to_LEFT_V6N017_2_0 ),
    .LEFT_V6S1(),
    .LEFT_V6S2(\net_do_reg[11]_LEFT_V6S2_to_LEFT_V6M214_2_0 ),
    .LEFT_V6S3(\net_do_reg[12]_LEFT_V6S3_to_LEFT_V6M314_2_0 ),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_16_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_16_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_16_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_16_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_16_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_16_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_16_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s1_w7.CONF = "0";
  defparam GSB_CNT_16_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_16_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_16_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(\net_do_reg[13]_W7_to_LEFT_E716_2_0 ),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(\net_do_reg[13]_N1_to_S116_3_0 ),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_16_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_16_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_16_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_16_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_16_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_16_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_16_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_16_2_0_inst.sps_o1.CONF = "110011110";
  defparam GSB_LFT_16_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_16_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_16_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_16_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_16_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_16_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_16_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_16_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_16_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_16_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_16_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_16_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_16_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_16_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_16_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_16_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_16_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_16_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_16_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(\net_do_reg[13]_W7_to_LEFT_E716_2_0 ),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_do_reg[13]_LEFT_O1_to_OUT16_2_0 ),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_13_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_13_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_13_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s14_w12.CONF = "0";
  defparam GSB_CNT_13_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s15_w17.CONF = "0";
  defparam GSB_CNT_13_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_13_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_do_reg[12]_W12_to_LEFT_E1213_2_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(\net_do_reg[11]_W17_to_LEFT_E1713_2_0 ),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(\net_do_reg[12]_N14_to_S1413_3_0 ),
    .S15(\net_do_reg[11]_N15_to_S1513_3_0 ),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_13_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_13_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_13_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_13_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_13_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_13_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_13_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_13_2_0_inst.sps_o2.CONF = "110100111";
  defparam GSB_LFT_13_2_0_inst.sps_o3.CONF = "110011011";
  defparam GSB_LFT_13_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_13_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_13_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(\net_do_reg[11]_W17_to_LEFT_E1713_2_0 ),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(\net_do_reg[12]_W12_to_LEFT_E1213_2_0 ),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(\net_do_reg[12]_LEFT_O2_to_OUT13_2_0 ),
    .LEFT_O3(\net_do_reg[11]_LEFT_O3_to_OUT13_2_0 ),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_5_14_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w2.CONF = "0000";
  defparam GSB_CNT_5_14_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_14_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_14_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s0.CONF = "0100";
  defparam GSB_CNT_5_14_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_14_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(\net_do_reg[11]_H6W2_to_H6E25_14_0 ),
    .H6E3(\net_do_reg[10]_H6W3_to_H6E35_14_0 ),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(\net_do_reg[11]_H6W2_to_H6E25_8_0 ),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(\net_do_reg[10]_V6S0_to_V6N011_14_0 ),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_h6w1.CONF = "0001";
  defparam GSB_CNT_5_8_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_h6w2.CONF = "0000";
  defparam GSB_CNT_5_8_0_inst.sps_h6w3.CONF = "0000";
  defparam GSB_CNT_5_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_8_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_8_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(\net_do_reg[11]_H6W2_to_H6E25_8_0 ),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_do_reg[5]_H6W1_to_H6M15_5_0 ),
    .H6W2(\net_do_reg[11]_H6W2_to_LEFT_H6E25_2_0 ),
    .H6W3(\net_do_reg[4]_H6W3_to_LEFT_H6E35_2_0 ),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[5]_LLH0_to_LLH05_8_0 ),
    .LLH6(\net_do_reg[4]_LLH6_to_LLH65_8_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_5_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_5_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_5_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_5_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_5_2_0_inst.sps_o3.CONF = "110101110";
  defparam GSB_LFT_5_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s2.CONF = "00111110";
  defparam GSB_LFT_5_2_0_inst.sps_v6s3.CONF = "00111110";
  defparam GSB_LFT_5_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_5_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_5_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(\net_do_reg[2]_W15_to_LEFT_E155_2_0 ),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(\net_do_reg[11]_H6W2_to_LEFT_H6E25_2_0 ),
    .LEFT_H6E3(\net_do_reg[4]_H6W3_to_LEFT_H6E35_2_0 ),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(\net_do_reg[11]_LEFT_V6S2_to_LEFT_V6N211_2_0 ),
    .LEFT_V6S3(\net_do_reg[4]_LEFT_V6S3_to_LEFT_V6M38_2_0 ),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(),
    .LEFT_O3(\net_do_reg[2]_LEFT_O3_to_OUT5_2_0 ),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_11_14_0_inst.sps_h6w0.CONF = "0100";
  defparam GSB_CNT_11_14_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_14_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_14_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_14_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_14_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_14_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_14_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_14_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_14_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(\net_do_reg[10]_H6W0_to_H6E011_8_0 ),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(\net_do_reg[10]_V6S0_to_V6N011_14_0 ),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_8_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s1.CONF = "0100";
  defparam GSB_CNT_11_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_8_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(\net_do_reg[10]_H6W0_to_H6E011_8_0 ),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(\net_do_reg[10]_V6S1_to_V6M114_8_0 ),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_14_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_h6w1.CONF = "0011";
  defparam GSB_CNT_14_8_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_14_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_14_8_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_14_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_14_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_14_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_14_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_14_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_14_8_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_do_reg[10]_H6W1_to_LEFT_H6E114_2_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_do_reg[10]_V6S1_to_V6M114_8_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_8_0_inst.sps_h6w0.CONF = "0001";
  defparam GSB_CNT_8_8_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w2.CONF = "0001";
  defparam GSB_CNT_8_8_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_8_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_8_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(\net_do_reg[8]_H6W0_to_LEFT_H6E08_2_0 ),
    .H6W1(),
    .H6W2(\net_do_reg[9]_H6W2_to_LEFT_H6E28_2_0 ),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[8]_LLH0_to_LLH08_8_0 ),
    .LLH6(\net_do_reg[9]_LLH6_to_LLH68_8_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_8_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_8_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_8_2_0_inst.sps_o1.CONF = "110110111";
  defparam GSB_LFT_8_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_8_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_8_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6s0.CONF = "00111110";
  defparam GSB_LFT_8_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6s2.CONF = "00111110";
  defparam GSB_LFT_8_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e12.CONF = "101";
  defparam GSB_LFT_8_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e22.CONF = "01";
  defparam GSB_LFT_8_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e3.CONF = "101";
  defparam GSB_LFT_8_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_8_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_8_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(\net_do_reg[4]_LEFT_E22_to_W228_3_0 ),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(\net_do_reg[9]_LEFT_E12_to_W128_3_0 ),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(\net_do_reg[8]_LEFT_E3_to_W38_3_0 ),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(\net_do_reg[8]_H6W0_to_LEFT_H6E08_2_0 ),
    .LEFT_H6E1(),
    .LEFT_H6E2(\net_do_reg[9]_H6W2_to_LEFT_H6E28_2_0 ),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(\net_do_reg[5]_H6W1_to_LEFT_H6M18_2_0 ),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(\net_do_reg[4]_LEFT_V6S3_to_LEFT_V6M38_2_0 ),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_do_reg[5]_LEFT_O1_to_OUT8_2_0 ),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_8_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s14_w12.CONF = "0";
  defparam GSB_CNT_8_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s20_w22.CONF = "0";
  defparam GSB_CNT_8_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s21_w3.CONF = "0";
  defparam GSB_CNT_8_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(\net_do_reg[8]_LEFT_E3_to_W38_3_0 ),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_do_reg[9]_LEFT_E12_to_W128_3_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(\net_do_reg[4]_LEFT_E22_to_W228_3_0 ),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(\net_do_reg[9]_S14_to_N149_3_0 ),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(\net_do_reg[4]_S20_to_N209_3_0 ),
    .S21(\net_do_reg[8]_S21_to_N219_3_0 ),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n14_w19.CONF = "0";
  defparam GSB_CNT_9_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n20_w1.CONF = "0";
  defparam GSB_CNT_9_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n21_w22.CONF = "0";
  defparam GSB_CNT_9_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s17_w23.CONF = "0";
  defparam GSB_CNT_9_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s2_w0.CONF = "0";
  defparam GSB_CNT_9_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(\net_do_reg[9]_S14_to_N149_3_0 ),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(\net_do_reg[4]_S20_to_N209_3_0 ),
    .N21(\net_do_reg[8]_S21_to_N219_3_0 ),
    .N22(),
    .N23(),
    .W0(\net_do_reg[7]_LEFT_E0_to_W09_3_0 ),
    .W1(\net_do_reg[4]_W1_to_LEFT_E19_2_0 ),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(\net_do_reg[9]_W19_to_LEFT_E199_2_0 ),
    .W20(),
    .W21(),
    .W22(\net_do_reg[8]_W22_to_LEFT_E229_2_0 ),
    .W23(\net_do_reg[6]_LEFT_E23_to_W239_3_0 ),
    .S0(),
    .S1(),
    .S2(\net_do_reg[7]_S2_to_N210_3_0 ),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(\net_do_reg[6]_S17_to_N1710_3_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_9_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_9_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_9_2_0_inst.sps_o1.CONF = "110101011";
  defparam GSB_LFT_9_2_0_inst.sps_o2.CONF = "110011110";
  defparam GSB_LFT_9_2_0_inst.sps_o3.CONF = "110001101";
  defparam GSB_LFT_9_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n3.CONF = "00111110";
  defparam GSB_LFT_9_2_0_inst.sps_v6s0.CONF = "00111110";
  defparam GSB_LFT_9_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_e0.CONF = "101";
  defparam GSB_LFT_9_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e23.CONF = "01";
  defparam GSB_LFT_9_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e0.CONF = "0111011";
  defparam GSB_LFT_9_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e2.CONF = "0111011";
  defparam GSB_LFT_9_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_9_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_9_2_0_inst (
    .LEFT_E23(\net_do_reg[6]_LEFT_E23_to_W239_3_0 ),
    .LEFT_E22(\net_do_reg[8]_W22_to_LEFT_E229_2_0 ),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(\net_do_reg[9]_W19_to_LEFT_E199_2_0 ),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(\net_do_reg[4]_W1_to_LEFT_E19_2_0 ),
    .LEFT_E0(\net_do_reg[7]_LEFT_E0_to_W09_3_0 ),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(\net_do_reg[7]_LLH6_to_LEFT_LLH09_2_0 ),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(\net_do_reg[6]_LLH0_to_LEFT_LLH69_2_0 ),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_do_reg[4]_LEFT_O1_to_OUT9_2_0 ),
    .LEFT_O2(\net_do_reg[9]_LEFT_O2_to_OUT9_2_0 ),
    .LEFT_O3(\net_do_reg[8]_LEFT_O3_to_OUT9_2_0 ),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_10_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n17_w18.CONF = "0";
  defparam GSB_CNT_10_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n2_w7.CONF = "0";
  defparam GSB_CNT_10_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(\net_do_reg[7]_S2_to_N210_3_0 ),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(\net_do_reg[6]_S17_to_N1710_3_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(\net_do_reg[7]_W7_to_LEFT_E710_2_0 ),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(\net_do_reg[6]_W18_to_LEFT_E1810_2_0 ),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_10_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_10_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_10_2_0_inst.sps_o1.CONF = "110011110";
  defparam GSB_LFT_10_2_0_inst.sps_o2.CONF = "110011101";
  defparam GSB_LFT_10_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_10_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_10_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_10_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(\net_do_reg[6]_W18_to_LEFT_E1810_2_0 ),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(\net_do_reg[7]_W7_to_LEFT_E710_2_0 ),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_do_reg[7]_LEFT_O1_to_OUT10_2_0 ),
    .LEFT_O2(\net_do_reg[6]_LEFT_O2_to_OUT10_2_0 ),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_5_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s1.CONF = "0011";
  defparam GSB_CNT_5_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_5_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(\net_do_reg[5]_H6W1_to_H6M15_5_0 ),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(\net_do_reg[5]_V6S1_to_V6M18_5_0 ),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w1.CONF = "0011";
  defparam GSB_CNT_8_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_5_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_do_reg[5]_H6W1_to_LEFT_H6M18_2_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_do_reg[5]_V6S1_to_V6M18_5_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_h6w1.CONF = "0001";
  defparam GSB_CNT_4_8_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_8_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_8_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_do_reg[3]_H6W1_to_LEFT_H6E14_2_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_do_reg[3]_LLH0_to_LLH04_8_0 ),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_4_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_4_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_4_2_0_inst.sps_o1.CONF = "110111110";
  defparam GSB_LFT_4_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_4_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_4_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n1.CONF = "00111110";
  defparam GSB_LFT_4_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e8.CONF = "01";
  defparam GSB_LFT_4_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e0.CONF = "0111011";
  defparam GSB_LFT_4_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_4_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_4_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(\net_do_reg[2]_LEFT_E8_to_W84_3_0 ),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(\net_do_reg[3]_H6W1_to_LEFT_H6E14_2_0 ),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(\net_do_reg[2]_LLH6_to_LEFT_LLH04_2_0 ),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_do_reg[3]_LEFT_O1_to_OUT4_2_0 ),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_4_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s10_w8.CONF = "0";
  defparam GSB_CNT_4_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(\net_do_reg[2]_LEFT_E8_to_W84_3_0 ),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(\net_do_reg[2]_S10_to_N105_3_0 ),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n10_w15.CONF = "0";
  defparam GSB_CNT_5_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(\net_do_reg[2]_S10_to_N105_3_0 ),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(\net_do_reg[2]_W15_to_LEFT_E155_2_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_6_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_6_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_6_2_0_inst.sps_o1.CONF = "110111110";
  defparam GSB_LFT_6_2_0_inst.sps_o2.CONF = "110111110";
  defparam GSB_LFT_6_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_6_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e1.CONF = "0111011";
  defparam GSB_LFT_6_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e2.CONF = "0111011";
  defparam GSB_LFT_6_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_6_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_6_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(\net_do_reg[1]_LLH6_to_LEFT_LLH06_2_0 ),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(\net_do_reg[0]_LLH0_to_LEFT_LLH66_2_0 ),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_do_reg[1]_LEFT_O1_to_OUT6_2_0 ),
    .LEFT_O2(\net_do_reg[0]_LEFT_O2_to_OUT6_2_0 ),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  GSB_CLKC GSB_CLKC_18_28_0_inst (
    .CLKC_GCLK0(),
    .CLKC_GCLK1(\net_IBuf-clkpad-clk_CLKB_GCLK1_to_CLKC_GCLK118_28_0 ),
    .CLKC_GCLK2(),
    .CLKC_GCLK3(),
    .CLKC_HGCLK0(),
    .CLKC_HGCLK1(),
    .CLKC_HGCLK2(),
    .CLKC_HGCLK3(),
    .CLKC_VGCLK0(),
    .CLKC_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK112_28_0 ),
    .CLKC_VGCLK2(),
    .CLKC_VGCLK3()
  );

  defparam GSB_CLKV_12_28_0_inst.spbu_gclk_bufl0.CONF = "1";
  defparam GSB_CLKV_12_28_0_inst.spbu_gclk_bufl1.CONF = "0";
  defparam GSB_CLKV_12_28_0_inst.spbu_gclk_bufl2.CONF = "1";
  defparam GSB_CLKV_12_28_0_inst.spbu_gclk_bufl3.CONF = "1";
  defparam GSB_CLKV_12_28_0_inst.spbu_gclk_bufr0.CONF = "1";
  defparam GSB_CLKV_12_28_0_inst.spbu_gclk_bufr1.CONF = "1";
  defparam GSB_CLKV_12_28_0_inst.spbu_gclk_bufr2.CONF = "1";
  defparam GSB_CLKV_12_28_0_inst.spbu_gclk_bufr3.CONF = "1";
  GSB_CLKV GSB_CLKV_12_28_0_inst (
    .CLKV_VGCLK0(),
    .CLKV_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK112_28_0 ),
    .CLKV_VGCLK2(),
    .CLKV_VGCLK3(),
    .CLKV_GCLK_BUFL0(),
    .CLKV_GCLK_BUFL1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK112_21_0 ),
    .CLKV_GCLK_BUFL2(),
    .CLKV_GCLK_BUFL3(),
    .CLKV_GCLK_BUFR0(),
    .CLKV_GCLK_BUFR1(),
    .CLKV_GCLK_BUFR2(),
    .CLKV_GCLK_BUFR3()
  );

  defparam GSB_CLKV_11_28_0_inst.spbu_gclk_bufl0.CONF = "1";
  defparam GSB_CLKV_11_28_0_inst.spbu_gclk_bufl1.CONF = "0";
  defparam GSB_CLKV_11_28_0_inst.spbu_gclk_bufl2.CONF = "1";
  defparam GSB_CLKV_11_28_0_inst.spbu_gclk_bufl3.CONF = "1";
  defparam GSB_CLKV_11_28_0_inst.spbu_gclk_bufr0.CONF = "1";
  defparam GSB_CLKV_11_28_0_inst.spbu_gclk_bufr1.CONF = "1";
  defparam GSB_CLKV_11_28_0_inst.spbu_gclk_bufr2.CONF = "1";
  defparam GSB_CLKV_11_28_0_inst.spbu_gclk_bufr3.CONF = "1";
  GSB_CLKV GSB_CLKV_11_28_0_inst (
    .CLKV_VGCLK0(),
    .CLKV_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK112_28_0 ),
    .CLKV_VGCLK2(),
    .CLKV_VGCLK3(),
    .CLKV_GCLK_BUFL0(),
    .CLKV_GCLK_BUFL1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK111_21_0 ),
    .CLKV_GCLK_BUFL2(),
    .CLKV_GCLK_BUFL3(),
    .CLKV_GCLK_BUFR0(),
    .CLKV_GCLK_BUFR1(),
    .CLKV_GCLK_BUFR2(),
    .CLKV_GCLK_BUFR3()
  );

  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufl0.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufl1.CONF = "0";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufl2.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufl3.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufr0.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufr1.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufr2.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufr3.CONF = "1";
  GSB_CLKV GSB_CLKV_5_28_0_inst (
    .CLKV_VGCLK0(),
    .CLKV_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK112_28_0 ),
    .CLKV_VGCLK2(),
    .CLKV_VGCLK3(),
    .CLKV_GCLK_BUFL0(),
    .CLKV_GCLK_BUFL1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK15_21_0 ),
    .CLKV_GCLK_BUFL2(),
    .CLKV_GCLK_BUFL3(),
    .CLKV_GCLK_BUFR0(),
    .CLKV_GCLK_BUFR1(),
    .CLKV_GCLK_BUFR2(),
    .CLKV_GCLK_BUFR3()
  );

  defparam GSB_CLKV_8_28_0_inst.spbu_gclk_bufl0.CONF = "1";
  defparam GSB_CLKV_8_28_0_inst.spbu_gclk_bufl1.CONF = "0";
  defparam GSB_CLKV_8_28_0_inst.spbu_gclk_bufl2.CONF = "1";
  defparam GSB_CLKV_8_28_0_inst.spbu_gclk_bufl3.CONF = "1";
  defparam GSB_CLKV_8_28_0_inst.spbu_gclk_bufr0.CONF = "1";
  defparam GSB_CLKV_8_28_0_inst.spbu_gclk_bufr1.CONF = "1";
  defparam GSB_CLKV_8_28_0_inst.spbu_gclk_bufr2.CONF = "1";
  defparam GSB_CLKV_8_28_0_inst.spbu_gclk_bufr3.CONF = "1";
  GSB_CLKV GSB_CLKV_8_28_0_inst (
    .CLKV_VGCLK0(),
    .CLKV_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK112_28_0 ),
    .CLKV_VGCLK2(),
    .CLKV_VGCLK3(),
    .CLKV_GCLK_BUFL0(),
    .CLKV_GCLK_BUFL1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK18_21_0 ),
    .CLKV_GCLK_BUFL2(),
    .CLKV_GCLK_BUFL3(),
    .CLKV_GCLK_BUFR0(),
    .CLKV_GCLK_BUFR1(),
    .CLKV_GCLK_BUFR2(),
    .CLKV_GCLK_BUFR3()
  );

  defparam GSB_CLKV_9_28_0_inst.spbu_gclk_bufl0.CONF = "1";
  defparam GSB_CLKV_9_28_0_inst.spbu_gclk_bufl1.CONF = "0";
  defparam GSB_CLKV_9_28_0_inst.spbu_gclk_bufl2.CONF = "1";
  defparam GSB_CLKV_9_28_0_inst.spbu_gclk_bufl3.CONF = "1";
  defparam GSB_CLKV_9_28_0_inst.spbu_gclk_bufr0.CONF = "1";
  defparam GSB_CLKV_9_28_0_inst.spbu_gclk_bufr1.CONF = "1";
  defparam GSB_CLKV_9_28_0_inst.spbu_gclk_bufr2.CONF = "1";
  defparam GSB_CLKV_9_28_0_inst.spbu_gclk_bufr3.CONF = "1";
  GSB_CLKV GSB_CLKV_9_28_0_inst (
    .CLKV_VGCLK0(),
    .CLKV_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK112_28_0 ),
    .CLKV_VGCLK2(),
    .CLKV_VGCLK3(),
    .CLKV_GCLK_BUFL0(),
    .CLKV_GCLK_BUFL1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK19_21_0 ),
    .CLKV_GCLK_BUFL2(),
    .CLKV_GCLK_BUFL3(),
    .CLKV_GCLK_BUFR0(),
    .CLKV_GCLK_BUFR1(),
    .CLKV_GCLK_BUFR2(),
    .CLKV_GCLK_BUFR3()
  );

  defparam GSB_CLKV_4_28_0_inst.spbu_gclk_bufl0.CONF = "1";
  defparam GSB_CLKV_4_28_0_inst.spbu_gclk_bufl1.CONF = "0";
  defparam GSB_CLKV_4_28_0_inst.spbu_gclk_bufl2.CONF = "1";
  defparam GSB_CLKV_4_28_0_inst.spbu_gclk_bufl3.CONF = "1";
  defparam GSB_CLKV_4_28_0_inst.spbu_gclk_bufr0.CONF = "1";
  defparam GSB_CLKV_4_28_0_inst.spbu_gclk_bufr1.CONF = "1";
  defparam GSB_CLKV_4_28_0_inst.spbu_gclk_bufr2.CONF = "1";
  defparam GSB_CLKV_4_28_0_inst.spbu_gclk_bufr3.CONF = "1";
  GSB_CLKV GSB_CLKV_4_28_0_inst (
    .CLKV_VGCLK0(),
    .CLKV_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK112_28_0 ),
    .CLKV_VGCLK2(),
    .CLKV_VGCLK3(),
    .CLKV_GCLK_BUFL0(),
    .CLKV_GCLK_BUFL1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK14_21_0 ),
    .CLKV_GCLK_BUFL2(),
    .CLKV_GCLK_BUFL3(),
    .CLKV_GCLK_BUFR0(),
    .CLKV_GCLK_BUFR1(),
    .CLKV_GCLK_BUFR2(),
    .CLKV_GCLK_BUFR3()
  );

  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufl0.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufl1.CONF = "0";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufl2.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufl3.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufr0.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufr1.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufr2.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufr3.CONF = "1";
  GSB_CLKV GSB_CLKV_6_28_0_inst (
    .CLKV_VGCLK0(),
    .CLKV_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK112_28_0 ),
    .CLKV_VGCLK2(),
    .CLKV_VGCLK3(),
    .CLKV_GCLK_BUFL0(),
    .CLKV_GCLK_BUFL1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK16_21_0 ),
    .CLKV_GCLK_BUFL2(),
    .CLKV_GCLK_BUFL3(),
    .CLKV_GCLK_BUFR0(),
    .CLKV_GCLK_BUFR1(),
    .CLKV_GCLK_BUFR2(),
    .CLKV_GCLK_BUFR3()
  );

  defparam GSB_RHT_5_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh2.CONF = "01";
  defparam GSB_RHT_5_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_5_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_5_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_5_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_5_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_5_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_5_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_5_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_5_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(\net_Buf-pad-rstn_RIGHT_LLH2_to_LLH05_18_0 ),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(),
    .RIGHT_LLV6(),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(),
    .RIGHT_I3(\net_Buf-pad-rstn_IN_to_RIGHT_I35_54_0 ),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_5_18_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_18_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_18_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e1.CONF = "0000";
  defparam GSB_CNT_5_18_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_18_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(\net_Buf-pad-rstn_H6E1_to_H6M15_21_0 ),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_Buf-pad-rstn_RIGHT_LLH2_to_LLH05_18_0 ),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );
endmodule
