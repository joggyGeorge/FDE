
module inverter ( clk, rstn, cs, rd, di, empty, wr, do, full );
  input [15:0] di;
  output [15:0] do;
  input clk, rstn, cs, empty, full;
  output rd, wr;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63;
  wire   [15:0] di_q;
  wire   [15:0] di_d;
  wire   [15:0] do_d;
  wire   [2:0] cur_state;
  wire   [2:0] nxt_state;

  DFFRHQ \cur_state_reg[0]  ( .D(nxt_state[0]), .CK(clk), .RN(rstn), .Q(
        cur_state[0]) );
  DFFRHQ \cur_state_reg[1]  ( .D(nxt_state[1]), .CK(clk), .RN(rstn), .Q(
        cur_state[1]) );
  DFFRHQ \cur_state_reg[2]  ( .D(nxt_state[2]), .CK(clk), .RN(rstn), .Q(
        cur_state[2]) );
  DFFRHQ \di_q_reg[15]  ( .D(di_d[15]), .CK(clk), .RN(rstn), .Q(di_q[15]) );
  DFFRHQ \do_q_reg[15]  ( .D(do_d[15]), .CK(clk), .RN(rstn), .Q(do[15]) );
  DFFRHQ \di_q_reg[14]  ( .D(di_d[14]), .CK(clk), .RN(rstn), .Q(di_q[14]) );
  DFFRHQ \do_q_reg[14]  ( .D(do_d[14]), .CK(clk), .RN(rstn), .Q(do[14]) );
  DFFRHQ \di_q_reg[13]  ( .D(di_d[13]), .CK(clk), .RN(rstn), .Q(di_q[13]) );
  DFFRHQ \do_q_reg[13]  ( .D(do_d[13]), .CK(clk), .RN(rstn), .Q(do[13]) );
  DFFRHQ \di_q_reg[12]  ( .D(di_d[12]), .CK(clk), .RN(rstn), .Q(di_q[12]) );
  DFFRHQ \do_q_reg[12]  ( .D(do_d[12]), .CK(clk), .RN(rstn), .Q(do[12]) );
  DFFRHQ \di_q_reg[11]  ( .D(di_d[11]), .CK(clk), .RN(rstn), .Q(di_q[11]) );
  DFFRHQ \do_q_reg[11]  ( .D(do_d[11]), .CK(clk), .RN(rstn), .Q(do[11]) );
  DFFRHQ \di_q_reg[10]  ( .D(di_d[10]), .CK(clk), .RN(rstn), .Q(di_q[10]) );
  DFFRHQ \do_q_reg[10]  ( .D(do_d[10]), .CK(clk), .RN(rstn), .Q(do[10]) );
  DFFRHQ \di_q_reg[9]  ( .D(di_d[9]), .CK(clk), .RN(rstn), .Q(di_q[9]) );
  DFFRHQ \do_q_reg[9]  ( .D(do_d[9]), .CK(clk), .RN(rstn), .Q(do[9]) );
  DFFRHQ \di_q_reg[8]  ( .D(di_d[8]), .CK(clk), .RN(rstn), .Q(di_q[8]) );
  DFFRHQ \do_q_reg[8]  ( .D(do_d[8]), .CK(clk), .RN(rstn), .Q(do[8]) );
  DFFRHQ \di_q_reg[7]  ( .D(di_d[7]), .CK(clk), .RN(rstn), .Q(di_q[7]) );
  DFFRHQ \do_q_reg[7]  ( .D(do_d[7]), .CK(clk), .RN(rstn), .Q(do[7]) );
  DFFRHQ \di_q_reg[6]  ( .D(di_d[6]), .CK(clk), .RN(rstn), .Q(di_q[6]) );
  DFFRHQ \do_q_reg[6]  ( .D(do_d[6]), .CK(clk), .RN(rstn), .Q(do[6]) );
  DFFRHQ \di_q_reg[5]  ( .D(di_d[5]), .CK(clk), .RN(rstn), .Q(di_q[5]) );
  DFFRHQ \do_q_reg[5]  ( .D(do_d[5]), .CK(clk), .RN(rstn), .Q(do[5]) );
  DFFRHQ \di_q_reg[4]  ( .D(di_d[4]), .CK(clk), .RN(rstn), .Q(di_q[4]) );
  DFFRHQ \do_q_reg[4]  ( .D(do_d[4]), .CK(clk), .RN(rstn), .Q(do[4]) );
  DFFRHQ \di_q_reg[3]  ( .D(di_d[3]), .CK(clk), .RN(rstn), .Q(di_q[3]) );
  DFFRHQ \do_q_reg[3]  ( .D(do_d[3]), .CK(clk), .RN(rstn), .Q(do[3]) );
  DFFRHQ \di_q_reg[2]  ( .D(di_d[2]), .CK(clk), .RN(rstn), .Q(di_q[2]) );
  DFFRHQ \do_q_reg[2]  ( .D(do_d[2]), .CK(clk), .RN(rstn), .Q(do[2]) );
  DFFRHQ \di_q_reg[1]  ( .D(di_d[1]), .CK(clk), .RN(rstn), .Q(di_q[1]) );
  DFFRHQ \do_q_reg[1]  ( .D(do_d[1]), .CK(clk), .RN(rstn), .Q(do[1]) );
  DFFRHQ \di_q_reg[0]  ( .D(di_d[0]), .CK(clk), .RN(rstn), .Q(di_q[0]) );
  DFFRHQ \do_q_reg[0]  ( .D(do_d[0]), .CK(clk), .RN(rstn), .Q(do[0]) );
  OR3 U72 ( .A(cur_state[2]), .B(cur_state[0]), .C(n42), .Y(n35) );
  INV U73 ( .A(n47), .Y(n36) );
  INV U74 ( .A(n36), .Y(n37) );
  INV U75 ( .A(n35), .Y(n38) );
  OR2 U76 ( .A(n39), .B(n40), .Y(nxt_state[2]) );
  MX2 U77 ( .A(cur_state[2]), .B(n41), .S0(cur_state[0]), .Y(n40) );
  NOR2 U78 ( .A(full), .B(n42), .Y(n41) );
  INV U79 ( .A(n43), .Y(nxt_state[1]) );
  NOR3B U80 ( .AN(n44), .B(rd), .C(n39), .Y(n43) );
  NOR3B U81 ( .AN(cur_state[0]), .B(cur_state[2]), .C(cur_state[1]), .Y(rd) );
  NAND2 U82 ( .A(n44), .B(n45), .Y(nxt_state[0]) );
  AOI211 U83 ( .A0(cur_state[0]), .A1(n39), .B0(wr), .C0(n46), .Y(n45) );
  NOR4B U84 ( .AN(cs), .B(cur_state[1]), .C(cur_state[0]), .D(empty), .Y(n46)
         );
  NOR3B U85 ( .AN(cur_state[2]), .B(cur_state[1]), .C(cur_state[0]), .Y(wr) );
  NOR2B U86 ( .AN(cur_state[2]), .B(n42), .Y(n39) );
  AOI21 U87 ( .A0(n37), .A1(full), .B0(n38), .Y(n44) );
  MX2 U88 ( .A(do[9]), .B(n48), .S0(n37), .Y(do_d[9]) );
  INV U89 ( .A(di_q[9]), .Y(n48) );
  MX2 U90 ( .A(do[8]), .B(n49), .S0(n37), .Y(do_d[8]) );
  INV U91 ( .A(di_q[8]), .Y(n49) );
  MX2 U92 ( .A(do[7]), .B(n50), .S0(n37), .Y(do_d[7]) );
  INV U93 ( .A(di_q[7]), .Y(n50) );
  MX2 U94 ( .A(do[6]), .B(n51), .S0(n37), .Y(do_d[6]) );
  INV U95 ( .A(di_q[6]), .Y(n51) );
  MX2 U96 ( .A(do[5]), .B(n52), .S0(n37), .Y(do_d[5]) );
  INV U97 ( .A(di_q[5]), .Y(n52) );
  MX2 U98 ( .A(do[4]), .B(n53), .S0(n37), .Y(do_d[4]) );
  INV U99 ( .A(di_q[4]), .Y(n53) );
  MX2 U100 ( .A(do[3]), .B(n54), .S0(n37), .Y(do_d[3]) );
  INV U101 ( .A(di_q[3]), .Y(n54) );
  MX2 U102 ( .A(do[2]), .B(n55), .S0(n37), .Y(do_d[2]) );
  INV U103 ( .A(di_q[2]), .Y(n55) );
  MX2 U104 ( .A(do[1]), .B(n56), .S0(n37), .Y(do_d[1]) );
  INV U105 ( .A(di_q[1]), .Y(n56) );
  MX2 U106 ( .A(do[15]), .B(n57), .S0(n37), .Y(do_d[15]) );
  INV U107 ( .A(di_q[15]), .Y(n57) );
  MX2 U108 ( .A(do[14]), .B(n58), .S0(n37), .Y(do_d[14]) );
  INV U109 ( .A(di_q[14]), .Y(n58) );
  MX2 U110 ( .A(do[13]), .B(n59), .S0(n37), .Y(do_d[13]) );
  INV U111 ( .A(di_q[13]), .Y(n59) );
  MX2 U112 ( .A(do[12]), .B(n60), .S0(n37), .Y(do_d[12]) );
  INV U113 ( .A(di_q[12]), .Y(n60) );
  MX2 U114 ( .A(do[11]), .B(n61), .S0(n37), .Y(do_d[11]) );
  INV U115 ( .A(di_q[11]), .Y(n61) );
  MX2 U116 ( .A(do[10]), .B(n62), .S0(n37), .Y(do_d[10]) );
  INV U117 ( .A(di_q[10]), .Y(n62) );
  MX2 U118 ( .A(do[0]), .B(n63), .S0(n37), .Y(do_d[0]) );
  NOR3B U119 ( .AN(cur_state[0]), .B(cur_state[2]), .C(n42), .Y(n47) );
  INV U120 ( .A(di_q[0]), .Y(n63) );
  MX2 U121 ( .A(di_q[9]), .B(di[9]), .S0(n38), .Y(di_d[9]) );
  MX2 U122 ( .A(di_q[8]), .B(di[8]), .S0(n38), .Y(di_d[8]) );
  MX2 U123 ( .A(di_q[7]), .B(di[7]), .S0(n38), .Y(di_d[7]) );
  MX2 U124 ( .A(di_q[6]), .B(di[6]), .S0(n38), .Y(di_d[6]) );
  MX2 U125 ( .A(di_q[5]), .B(di[5]), .S0(n38), .Y(di_d[5]) );
  MX2 U126 ( .A(di_q[4]), .B(di[4]), .S0(n38), .Y(di_d[4]) );
  MX2 U127 ( .A(di_q[3]), .B(di[3]), .S0(n38), .Y(di_d[3]) );
  MX2 U128 ( .A(di_q[2]), .B(di[2]), .S0(n38), .Y(di_d[2]) );
  MX2 U129 ( .A(di_q[1]), .B(di[1]), .S0(n38), .Y(di_d[1]) );
  MX2 U130 ( .A(di_q[15]), .B(di[15]), .S0(n38), .Y(di_d[15]) );
  MX2 U131 ( .A(di_q[14]), .B(di[14]), .S0(n38), .Y(di_d[14]) );
  MX2 U132 ( .A(di_q[13]), .B(di[13]), .S0(n38), .Y(di_d[13]) );
  MX2 U133 ( .A(di_q[12]), .B(di[12]), .S0(n38), .Y(di_d[12]) );
  MX2 U134 ( .A(di_q[11]), .B(di[11]), .S0(n38), .Y(di_d[11]) );
  MX2 U135 ( .A(di_q[10]), .B(di[10]), .S0(n38), .Y(di_d[10]) );
  MX2 U136 ( .A(di_q[0]), .B(di[0]), .S0(n38), .Y(di_d[0]) );
  INV U137 ( .A(cur_state[1]), .Y(n42) );
endmodule

