//-------------------------------------------------------------------
//
//  COPYRIGHT (C) 2012, Renfeng Dou, Fudan University
//
//  THIS FILE MAY NOT BE MODIFIED OR REDISTRIBUTED WITHOUT THE
//  EXPRESSED WRITTEN CONSENT OF Renfeng Dou
//
//  Renfeng Dou			    email:12212020002@fudan.edu.cn
//  Fudan University          www.fudan.edu.cn
//-------------------------------------------------------------------
// Filename       : left_pic_rom.v
// Author         : Renfeng Dou
// Created        : 2012/10/25 0:00:00
// Description    : ROM file for VeriInstrument Graphic LCD
//
//-------------------------------------------------------------------

//synopsys_translate_off
`timescale 1ns/1ns
//synopsys_translate_on

module left_pic_rom(
                  clk,
                  rst_n,
                  sync_i,
                  en_i,
                  d_o,
                  length_o
);

input         clk;
input         rst_n;
input         sync_i;
input         en_i;
output [8:0]  d_o;
output [9:0]  length_o;

reg [9:0]     counter_r;

reg [8:0]     d_o;
reg [9:0]     length_o;

always @ (counter_r)
begin
  case(counter_r)
  10'd0: d_o =   {8'h3e,1'b0};
  10'd1: d_o =   {8'hb9,1'b0};
  10'd2: d_o =   {8'h4f,1'b0};
  10'd3: d_o =   {8'h01,1'b1};
  10'd4: d_o =   {8'h03,1'b1};
  10'd5: d_o =   {8'h06,1'b1};
  10'd6: d_o =   {8'h0e,1'b1};
  10'd7: d_o =   {8'h08,1'b1};
  10'd8: d_o =   {8'h18,1'b1};
  10'd9: d_o =   {8'h30,1'b1};
  10'd10: d_o =   {8'h37,1'b1};
  10'd11: d_o =   {8'h32,1'b1};
  10'd12: d_o =   {8'h61,1'b1};
  10'd13: d_o =   {8'h46,1'b1};
  10'd14: d_o =   {8'h4e,1'b1};
  10'd15: d_o =   {8'h51,1'b1};
  10'd16: d_o =   {8'hd0,1'b1};
  10'd17: d_o =   {8'hf8,1'b1};
  10'd18: d_o =   {8'hc3,1'b1};
  10'd19: d_o =   {8'hbc,1'b1};
  10'd20: d_o =   {8'h81,1'b1};
  10'd21: d_o =   {8'h81,1'b1};
  10'd22: d_o =   {8'h81,1'b1};
  10'd23: d_o =   {8'hbc,1'b1};
  10'd24: d_o =   {8'ha0,1'b1};
  10'd25: d_o =   {8'hf4,1'b1};
  10'd26: d_o =   {8'h55,1'b1};
  10'd27: d_o =   {8'h5f,1'b1};
  10'd28: d_o =   {8'h40,1'b1};
  10'd29: d_o =   {8'h60,1'b1};
  10'd30: d_o =   {8'h60,1'b1};
  10'd31: d_o =   {8'h30,1'b1};
  10'd32: d_o =   {8'h30,1'b1};
  10'd33: d_o =   {8'h30,1'b1};
  10'd34: d_o =   {8'h08,1'b1};
  10'd35: d_o =   {8'h0c,1'b1};
  10'd36: d_o =   {8'h06,1'b1};
  10'd37: d_o =   {8'h06,1'b1};
  10'd38: d_o =   {8'h01,1'b1};
  10'd39: d_o =   {8'hba,1'b0};
  10'd40: d_o =   {8'h49,1'b0};
  10'd41: d_o =   {8'h01,1'b1};
  10'd42: d_o =   {8'h03,1'b1};
  10'd43: d_o =   {8'h0e,1'b1};
  10'd44: d_o =   {8'h39,1'b1};
  10'd45: d_o =   {8'h30,1'b1};
  10'd46: d_o =   {8'hc0,1'b1};
  10'd47: d_o =   {8'h90,1'b1};
  10'd48: d_o =   {8'h08,1'b1};
  10'd49: d_o =   {8'h00,1'b1};
  10'd50: d_o =   {8'h7c,1'b1};
  10'd51: d_o =   {8'h21,1'b1};
  10'd52: d_o =   {8'h21,1'b1};
  10'd53: d_o =   {8'h16,1'b1};
  10'd54: d_o =   {8'he4,1'b1};
  10'd55: d_o =   {8'h28,1'b1};
  10'd56: d_o =   {8'h18,1'b1};
  10'd57: d_o =   {8'h97,1'b1};
  10'd58: d_o =   {8'haf,1'b1};
  10'd59: d_o =   {8'h3c,1'b1};
  10'd60: d_o =   {8'h38,1'b1};
  10'd61: d_o =   {8'h58,1'b1};
  10'd62: d_o =   {8'h5f,1'b1};
  10'd63: d_o =   {8'h5f,1'b1};
  10'd64: d_o =   {8'hd8,1'b1};
  10'd65: d_o =   {8'hd8,1'b1};
  10'd66: d_o =   {8'h5e,1'b1};
  10'd67: d_o =   {8'h4f,1'b1};
  10'd68: d_o =   {8'h47,1'b1};
  10'd69: d_o =   {8'h40,1'b1};
  10'd70: d_o =   {8'h27,1'b1};
  10'd71: d_o =   {8'hbf,1'b1};
  10'd72: d_o =   {8'h3f,1'b1};
  10'd73: d_o =   {8'h10,1'b1};
  10'd74: d_o =   {8'h18,1'b1};
  10'd75: d_o =   {8'h08,1'b1};
  10'd76: d_o =   {8'h04,1'b1};
  10'd77: d_o =   {8'h02,1'b1};
  10'd78: d_o =   {8'h01,1'b1};
  10'd79: d_o =   {8'h00,1'b1};
  10'd80: d_o =   {8'h02,1'b1};
  10'd81: d_o =   {8'h02,1'b1};
  10'd82: d_o =   {8'h04,1'b1};
  10'd83: d_o =   {8'hcc,1'b1};
  10'd84: d_o =   {8'hc8,1'b1};
  10'd85: d_o =   {8'h30,1'b1};
  10'd86: d_o =   {8'h1c,1'b1};
  10'd87: d_o =   {8'h06,1'b1};
  10'd88: d_o =   {8'h03,1'b1};
  10'd89: d_o =   {8'hbb,1'b0};
  10'd90: d_o =   {8'h48,1'b0};
  10'd91: d_o =   {8'h3f,1'b1};
  10'd92: d_o =   {8'hf0,1'b1};
  10'd93: d_o =   {8'hc0,1'b1};
  10'd94: d_o =   {8'h11,1'b1};
  10'd95: d_o =   {8'h80,1'b1};
  10'd96: d_o =   {8'h88,1'b1};
  10'd97: d_o =   {8'h08,1'b1};
  10'd98: d_o =   {8'h4b,1'b1};
  10'd99: d_o =   {8'h21,1'b1};
  10'd100: d_o =   {8'h0f,1'b1};
  10'd101: d_o =   {8'h70,1'b1};
  10'd102: d_o =   {8'h80,1'b1};
  10'd103: d_o =   {8'h80,1'b1};
  10'd104: d_o =   {8'h01,1'b1};
  10'd105: d_o =   {8'h03,1'b1};
  10'd106: d_o =   {8'h03,1'b1};
  10'd107: d_o =   {8'h06,1'b1};
  10'd108: d_o =   {8'hf0,1'b1};
  10'd109: d_o =   {8'hf0,1'b1};
  10'd110: d_o =   {8'h31,1'b1};
  10'd111: d_o =   {8'h3f,1'b1};
  10'd112: d_o =   {8'h3f,1'b1};
  10'd113: d_o =   {8'hfe,1'b1};
  10'd114: d_o =   {8'hf8,1'b1};
  10'd115: d_o =   {8'h39,1'b1};
  10'd116: d_o =   {8'h39,1'b1};
  10'd117: d_o =   {8'hf9,1'b1};
  10'd118: d_o =   {8'hf1,1'b1};
  10'd119: d_o =   {8'hf1,1'b1};
  10'd120: d_o =   {8'h03,1'b1};
  10'd121: d_o =   {8'hff,1'b1};
  10'd122: d_o =   {8'hff,1'b1};
  10'd123: d_o =   {8'hc3,1'b1};
  10'd124: d_o =   {8'h01,1'b1};
  10'd125: d_o =   {8'h01,1'b1};
  10'd126: d_o =   {8'h01,1'b1};
  10'd127: d_o =   {8'h01,1'b1};
  10'd128: d_o =   {8'h01,1'b1};
  10'd129: d_o =   {8'h81,1'b1};
  10'd130: d_o =   {8'h40,1'b1};
  10'd131: d_o =   {8'h1c,1'b1};
  10'd132: d_o =   {8'h07,1'b1};
  10'd133: d_o =   {8'h08,1'b1};
  10'd134: d_o =   {8'h12,1'b1};
  10'd135: d_o =   {8'h32,1'b1};
  10'd136: d_o =   {8'h02,1'b1};
  10'd137: d_o =   {8'h04,1'b1};
  10'd138: d_o =   {8'h18,1'b1};
  10'd139: d_o =   {8'hc0,1'b1};
  10'd140: d_o =   {8'h7f,1'b1};
  10'd141: d_o =   {8'h0f,1'b1};
  10'd142: d_o =   {8'hbc,1'b0};
  10'd143: d_o =   {8'h48,1'b0};
  10'd144: d_o =   {8'hff,1'b1};
  10'd145: d_o =   {8'h01,1'b1};
  10'd146: d_o =   {8'h20,1'b1};
  10'd147: d_o =   {8'h25,1'b1};
  10'd148: d_o =   {8'ha4,1'b1};
  10'd149: d_o =   {8'he4,1'b1};
  10'd150: d_o =   {8'h24,1'b1};
  10'd151: d_o =   {8'h0c,1'b1};
  10'd152: d_o =   {8'hf0,1'b1};
  10'd153: d_o =   {8'hfe,1'b1};
  10'd154: d_o =   {8'h41,1'b1};
  10'd155: d_o =   {8'hc0,1'b1};
  10'd156: d_o =   {8'hc0,1'b1};
  10'd157: d_o =   {8'hc0,1'b1};
  10'd158: d_o =   {8'hff,1'b1};
  10'd159: d_o =   {8'hff,1'b1};
  10'd160: d_o =   {8'hc7,1'b1};
  10'd161: d_o =   {8'hdf,1'b1};
  10'd162: d_o =   {8'hd8,1'b1};
  10'd163: d_o =   {8'hff,1'b1};
  10'd164: d_o =   {8'he7,1'b1};
  10'd165: d_o =   {8'hc0,1'b1};
  10'd166: d_o =   {8'hcf,1'b1};
  10'd167: d_o =   {8'hd8,1'b1};
  10'd168: d_o =   {8'hdc,1'b1};
  10'd169: d_o =   {8'hdf,1'b1};
  10'd170: d_o =   {8'hc0,1'b1};
  10'd171: d_o =   {8'h87,1'b1};
  10'd172: d_o =   {8'h8f,1'b1};
  10'd173: d_o =   {8'h83,1'b1};
  10'd174: d_o =   {8'hbf,1'b1};
  10'd175: d_o =   {8'hbf,1'b1};
  10'd176: d_o =   {8'h83,1'b1};
  10'd177: d_o =   {8'h9f,1'b1};
  10'd178: d_o =   {8'hbd,1'b1};
  10'd179: d_o =   {8'h81,1'b1};
  10'd180: d_o =   {8'h80,1'b1};
  10'd181: d_o =   {8'hc0,1'b1};
  10'd182: d_o =   {8'hc0,1'b1};
  10'd183: d_o =   {8'hc0,1'b1};
  10'd184: d_o =   {8'h07,1'b1};
  10'd185: d_o =   {8'hfc,1'b1};
  10'd186: d_o =   {8'h00,1'b1};
  10'd187: d_o =   {8'h0a,1'b1};
  10'd188: d_o =   {8'h1a,1'b1};
  10'd189: d_o =   {8'h19,1'b1};
  10'd190: d_o =   {8'h09,1'b1};
  10'd191: d_o =   {8'h08,1'b1};
  10'd192: d_o =   {8'h00,1'b1};
  10'd193: d_o =   {8'hff,1'b1};
  10'd194: d_o =   {8'hfe,1'b1};
  10'd195: d_o =   {8'hbd,1'b0};
  10'd196: d_o =   {8'h49,1'b0};
  10'd197: d_o =   {8'hf0,1'b1};
  10'd198: d_o =   {8'h78,1'b1};
  10'd199: d_o =   {8'h8e,1'b1};
  10'd200: d_o =   {8'h83,1'b1};
  10'd201: d_o =   {8'h89,1'b1};
  10'd202: d_o =   {8'ha6,1'b1};
  10'd203: d_o =   {8'hc4,1'b1};
  10'd204: d_o =   {8'h8c,1'b1};
  10'd205: d_o =   {8'h0a,1'b1};
  10'd206: d_o =   {8'h80,1'b1};
  10'd207: d_o =   {8'h66,1'b1};
  10'd208: d_o =   {8'h31,1'b1};
  10'd209: d_o =   {8'h09,1'b1};
  10'd210: d_o =   {8'hfc,1'b1};
  10'd211: d_o =   {8'hf6,1'b1};
  10'd212: d_o =   {8'hf1,1'b1};
  10'd213: d_o =   {8'hf9,1'b1};
  10'd214: d_o =   {8'h19,1'b1};
  10'd215: d_o =   {8'hf8,1'b1};
  10'd216: d_o =   {8'hf0,1'b1};
  10'd217: d_o =   {8'h00,1'b1};
  10'd218: d_o =   {8'hf8,1'b1};
  10'd219: d_o =   {8'h18,1'b1};
  10'd220: d_o =   {8'h78,1'b1};
  10'd221: d_o =   {8'hf8,1'b1};
  10'd222: d_o =   {8'h00,1'b1};
  10'd223: d_o =   {8'hc8,1'b1};
  10'd224: d_o =   {8'hd8,1'b1};
  10'd225: d_o =   {8'hf8,1'b1};
  10'd226: d_o =   {8'hd8,1'b1};
  10'd227: d_o =   {8'h98,1'b1};
  10'd228: d_o =   {8'hf9,1'b1};
  10'd229: d_o =   {8'hc1,1'b1};
  10'd230: d_o =   {8'hc1,1'b1};
  10'd231: d_o =   {8'hc6,1'b1};
  10'd232: d_o =   {8'h48,1'b1};
  10'd233: d_o =   {8'h48,1'b1};
  10'd234: d_o =   {8'h30,1'b1};
  10'd235: d_o =   {8'hc8,1'b1};
  10'd236: d_o =   {8'h10,1'b1};
  10'd237: d_o =   {8'h0e,1'b1};
  10'd238: d_o =   {8'h01,1'b1};
  10'd239: d_o =   {8'h01,1'b1};
  10'd240: d_o =   {8'h00,1'b1};
  10'd241: d_o =   {8'h01,1'b1};
  10'd242: d_o =   {8'h06,1'b1};
  10'd243: d_o =   {8'h0e,1'b1};
  10'd244: d_o =   {8'h70,1'b1};
  10'd245: d_o =   {8'h80,1'b1};
  10'd246: d_o =   {8'hbe,1'b0};
  10'd247: d_o =   {8'h4d,1'b0};
  10'd248: d_o =   {8'hc0,1'b1};
  10'd249: d_o =   {8'he0,1'b1};
  10'd250: d_o =   {8'h30,1'b1};
  10'd251: d_o =   {8'h18,1'b1};
  10'd252: d_o =   {8'h1c,1'b1};
  10'd253: d_o =   {8'h24,1'b1};
  10'd254: d_o =   {8'hd2,1'b1};
  10'd255: d_o =   {8'hd2,1'b1};
  10'd256: d_o =   {8'h63,1'b1};
  10'd257: d_o =   {8'hc1,1'b1};
  10'd258: d_o =   {8'hc1,1'b1};
  10'd259: d_o =   {8'h06,1'b1};
  10'd260: d_o =   {8'h08,1'b1};
  10'd261: d_o =   {8'h0a,1'b1};
  10'd262: d_o =   {8'hb8,1'b1};
  10'd263: d_o =   {8'hc1,1'b1};
  10'd264: d_o =   {8'hdf,1'b1};
  10'd265: d_o =   {8'h40,1'b1};
  10'd266: d_o =   {8'h41,1'b1};
  10'd267: d_o =   {8'h5f,1'b1};
  10'd268: d_o =   {8'h5d,1'b1};
  10'd269: d_o =   {8'h41,1'b1};
  10'd270: d_o =   {8'h40,1'b1};
  10'd271: d_o =   {8'h41,1'b1};
  10'd272: d_o =   {8'hff,1'b1};
  10'd273: d_o =   {8'h84,1'b1};
  10'd274: d_o =   {8'h80,1'b1};
  10'd275: d_o =   {8'h02,1'b1};
  10'd276: d_o =   {8'h00,1'b1};
  10'd277: d_o =   {8'h00,1'b1};
  10'd278: d_o =   {8'h01,1'b1};
  10'd279: d_o =   {8'h01,1'b1};
  10'd280: d_o =   {8'h03,1'b1};
  10'd281: d_o =   {8'h02,1'b1};
  10'd282: d_o =   {8'h04,1'b1};
  10'd283: d_o =   {8'h0c,1'b1};
  10'd284: d_o =   {8'h18,1'b1};
  10'd285: d_o =   {8'h10,1'b1};
  10'd286: d_o =   {8'h60,1'b1};
  10'd287: d_o =   {8'hc0,1'b1};
  10'd288: d_o =   {8'h80,1'b1};
  10'd289: d_o =   {8'hbf,1'b0};
  10'd290: d_o =   {8'h56,1'b0};
  10'd291: d_o =   {8'h80,1'b1};
  10'd292: d_o =   {8'h80,1'b1};
  10'd293: d_o =   {8'h80,1'b1};
  10'd294: d_o =   {8'hc0,1'b1};
  10'd295: d_o =   {8'h40,1'b1};
  10'd296: d_o =   {8'h40,1'b1};
  10'd297: d_o =   {8'h40,1'b1};
  10'd298: d_o =   {8'h40,1'b1};
  10'd299: d_o =   {8'h40,1'b1};
  10'd300: d_o =   {8'h60,1'b1};
  10'd301: d_o =   {8'h20,1'b1};
  10'd302: d_o =   {8'h20,1'b1};
  10'd303: d_o =   {8'h60,1'b1};
  10'd304: d_o =   {8'h60,1'b1};
  10'd305: d_o =   {8'h40,1'b1};
  10'd306: d_o =   {8'h40,1'b1};
  10'd307: d_o =   {8'h40,1'b1};
  10'd308: d_o =   {8'h40,1'b1};
  10'd309: d_o =   {8'h40,1'b1};
  10'd310: d_o =   {8'hc0,1'b1};
  10'd311: d_o =   {8'h80,1'b1};
  10'd312: d_o =   {8'h80,1'b1};
  10'd313: d_o =   {8'h3f,1'b0};
  default:d_o =   {8'h00,1'b1};
  endcase
end

always @ (posedge clk or negedge rst_n)
begin
  if(!rst_n)
      begin
          length_o    <= 10'd313;
          counter_r   <= 10'd0;
      end
  else
      begin                         // sync = 0 & en_i = 0 then couter++
          length_o  <= 10'd313;
          if(sync_i)
              counter_r   <= 10'd0;
          else if(!en_i)
              if(counter_r<length_o)
                  counter_r   <= counter_r + 1'b1;
      end
end

endmodule
