
module top ( clk, rst_n, auto_i, manual_i, graphic_lcd_d, graphic_lcd_rw, 
        graphic_lcd_en, graphic_lcd_di, graphic_lcd_rst, graphic_lcd_cs1, 
        graphic_lcd_cs2 );
  output [7:0] graphic_lcd_d;
  input clk, rst_n, auto_i, manual_i;
  output graphic_lcd_rw, graphic_lcd_en, graphic_lcd_di, graphic_lcd_rst,
         graphic_lcd_cs1, graphic_lcd_cs2;
  wire   sync_right, mode, _0_net_, refresh, \g_l_d1/counter[0] ,
         \g_l_d1/counter[1] , \g_l_d1/counter[2] , \g_l_d1/counter[3] ,
         \g_l_d1/counter[4] , \g_l_d1/counter[5] , \g_l_d1/counter[6] ,
         \g_l_d1/counter[7] , \g_l_d1/counter[8] , \g_l_d1/counter[9] ,
         \g_l_d1/state[0] , \g_l_d1/state[1] , \g_l_d1/state[2] ,
         \g_l_d1/*Logic0* , \l_p_r/N2857 , \l_p_r/N2856 , \l_p_r/N2855 ,
         \l_p_r/N2854 , \l_p_r/N2853 , \l_p_r/N2852 , \l_p_r/N2851 ,
         \l_p_r/N2850 , \l_p_r/N2849 , \l_p_r/counter_r[0] ,
         \l_p_r/counter_r[1] , \l_p_r/counter_r[2] , \l_p_r/counter_r[3] ,
         \l_p_r/counter_r[4] , \l_p_r/counter_r[5] , \l_p_r/counter_r[6] ,
         \l_p_r/counter_r[7] , \l_p_r/counter_r[8] , \r_p_r/N3466 ,
         \r_p_r/N3465 , \r_p_r/N3464 , \r_p_r/N3463 , \r_p_r/N3462 ,
         \r_p_r/N3461 , \r_p_r/N3460 , \r_p_r/N3459 , \r_p_r/N3458 ,
         \r_p_r/counter_r[0] , \r_p_r/counter_r[1] , \r_p_r/counter_r[2] ,
         \r_p_r/counter_r[3] , \r_p_r/counter_r[4] , \r_p_r/counter_r[5] ,
         \r_p_r/counter_r[6] , \r_p_r/counter_r[7] , \r_p_r/counter_r[8] ,
         \re_detect1/sample_r[0] , \re_detect1/sample_r[1] , n86, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n208, n209, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n227, n228, n230, n231, n232,
         n233, n234, n235, n236, n237, n239, n240, n241, n242, n243, n244,
         n245, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n359, n360, n361, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n649, n651, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411;
  wire   [13:0] \clk_div1/counter ;
  assign graphic_lcd_rw = \g_l_d1/*Logic0* ;

  DFFRHQ \clk_div1/counter_reg[14]  ( .D(n1341), .CK(clk), .RN(rst_n), .Q(
        refresh) );
  DFFRHQ \clk_div1/counter_reg[0]  ( .D(n1355), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [0]) );
  DFFRHQ \clk_div1/counter_reg[1]  ( .D(n1354), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [1]) );
  DFFRHQ \clk_div1/counter_reg[2]  ( .D(n1353), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [2]) );
  DFFRHQ \clk_div1/counter_reg[3]  ( .D(n1352), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [3]) );
  DFFRHQ \clk_div1/counter_reg[4]  ( .D(n1351), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [4]) );
  DFFRHQ \clk_div1/counter_reg[5]  ( .D(n1350), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [5]) );
  DFFRHQ \clk_div1/counter_reg[6]  ( .D(n1349), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [6]) );
  DFFRHQ \clk_div1/counter_reg[7]  ( .D(n1348), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [7]) );
  DFFRHQ \clk_div1/counter_reg[8]  ( .D(n1347), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [8]) );
  DFFRHQ \clk_div1/counter_reg[9]  ( .D(n1346), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [9]) );
  DFFRHQ \clk_div1/counter_reg[10]  ( .D(n1345), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [10]) );
  DFFRHQ \clk_div1/counter_reg[11]  ( .D(n1344), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [11]) );
  DFFRHQ \clk_div1/counter_reg[12]  ( .D(n1343), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [12]) );
  DFFRHQ \clk_div1/counter_reg[13]  ( .D(n1342), .CK(clk), .RN(rst_n), .Q(
        \clk_div1/counter [13]) );
  DFFRHQ \re_detect1/sample_r_reg[0]  ( .D(_0_net_), .CK(clk), .RN(rst_n), .Q(
        \re_detect1/sample_r[0] ) );
  DFFRHQ \re_detect1/sample_r_reg[1]  ( .D(\re_detect1/sample_r[0] ), .CK(clk), 
        .RN(rst_n), .Q(\re_detect1/sample_r[1] ) );
  DFFRHQ \g_l_d1/state_reg[1]  ( .D(n205), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/state[1] ) );
  DFFRHQ \g_l_d1/state_reg[0]  ( .D(n201), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/state[0] ) );
  DFFRHQ \g_l_d1/counter_reg[9]  ( .D(n203), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/counter[9] ) );
  DFFRHQ \g_l_d1/state_reg[2]  ( .D(n202), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/state[2] ) );
  DFFSHQ \g_l_d1/lcd_rst_o_reg  ( .D(n190), .CK(clk), .SN(rst_n), .Q(
        graphic_lcd_rst) );
  DFFRHQ \g_l_d1/cs1_reg  ( .D(n191), .CK(clk), .RN(rst_n), .Q(graphic_lcd_cs1) );
  DFFRHQ \g_l_d1/sync_right_reg  ( .D(n206), .CK(clk), .RN(rst_n), .Q(
        sync_right) );
  DFFRHQ \g_l_d1/lcd_en_o_reg  ( .D(n204), .CK(clk), .RN(rst_n), .Q(
        graphic_lcd_en) );
  DFFRHQ \g_l_d1/counter_reg[0]  ( .D(n192), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/counter[0] ) );
  DFFRHQ \g_l_d1/counter_reg[1]  ( .D(n193), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/counter[1] ) );
  DFFRHQ \g_l_d1/counter_reg[2]  ( .D(n194), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/counter[2] ) );
  DFFRHQ \g_l_d1/counter_reg[3]  ( .D(n195), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/counter[3] ) );
  DFFRHQ \g_l_d1/counter_reg[4]  ( .D(n196), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/counter[4] ) );
  DFFRHQ \g_l_d1/counter_reg[5]  ( .D(n197), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/counter[5] ) );
  DFFRHQ \g_l_d1/counter_reg[6]  ( .D(n198), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/counter[6] ) );
  DFFRHQ \g_l_d1/counter_reg[7]  ( .D(n199), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/counter[7] ) );
  DFFRHQ \g_l_d1/counter_reg[8]  ( .D(n200), .CK(clk), .RN(rst_n), .Q(
        \g_l_d1/counter[8] ) );
  DFFRHQ \g_l_d1/mode_reg  ( .D(n86), .CK(clk), .RN(rst_n), .Q(mode) );
  DFFRHQ \r_p_r/counter_r_reg[0]  ( .D(n178), .CK(clk), .RN(rst_n), .Q(
        \r_p_r/counter_r[0] ) );
  DFFRHQ \r_p_r/counter_r_reg[1]  ( .D(n177), .CK(clk), .RN(rst_n), .Q(
        \r_p_r/counter_r[1] ) );
  DFFRHQ \r_p_r/counter_r_reg[2]  ( .D(n176), .CK(clk), .RN(rst_n), .Q(
        \r_p_r/counter_r[2] ) );
  DFFRHQ \r_p_r/counter_r_reg[3]  ( .D(n175), .CK(clk), .RN(rst_n), .Q(
        \r_p_r/counter_r[3] ) );
  DFFRHQ \r_p_r/counter_r_reg[4]  ( .D(n174), .CK(clk), .RN(rst_n), .Q(
        \r_p_r/counter_r[4] ) );
  DFFRHQ \r_p_r/counter_r_reg[5]  ( .D(n173), .CK(clk), .RN(rst_n), .Q(
        \r_p_r/counter_r[5] ) );
  DFFRHQ \r_p_r/counter_r_reg[6]  ( .D(n172), .CK(clk), .RN(rst_n), .Q(
        \r_p_r/counter_r[6] ) );
  DFFRHQ \r_p_r/counter_r_reg[7]  ( .D(n171), .CK(clk), .RN(rst_n), .Q(
        \r_p_r/counter_r[7] ) );
  DFFRHQ \r_p_r/counter_r_reg[8]  ( .D(n170), .CK(clk), .RN(rst_n), .Q(
        \r_p_r/counter_r[8] ) );
  DFFRHQ \l_p_r/counter_r_reg[0]  ( .D(n188), .CK(clk), .RN(rst_n), .Q(
        \l_p_r/counter_r[0] ) );
  DFFRHQ \l_p_r/counter_r_reg[1]  ( .D(n187), .CK(clk), .RN(rst_n), .Q(
        \l_p_r/counter_r[1] ) );
  DFFRHQ \l_p_r/counter_r_reg[2]  ( .D(n186), .CK(clk), .RN(rst_n), .Q(
        \l_p_r/counter_r[2] ) );
  DFFRHQ \l_p_r/counter_r_reg[3]  ( .D(n185), .CK(clk), .RN(rst_n), .Q(
        \l_p_r/counter_r[3] ) );
  DFFRHQ \l_p_r/counter_r_reg[4]  ( .D(n184), .CK(clk), .RN(rst_n), .Q(
        \l_p_r/counter_r[4] ) );
  DFFRHQ \l_p_r/counter_r_reg[5]  ( .D(n183), .CK(clk), .RN(rst_n), .Q(
        \l_p_r/counter_r[5] ) );
  DFFRHQ \l_p_r/counter_r_reg[6]  ( .D(n182), .CK(clk), .RN(rst_n), .Q(
        \l_p_r/counter_r[6] ) );
  DFFRHQ \l_p_r/counter_r_reg[7]  ( .D(n181), .CK(clk), .RN(rst_n), .Q(
        \l_p_r/counter_r[7] ) );
  DFFRHQ \l_p_r/counter_r_reg[8]  ( .D(n180), .CK(clk), .RN(rst_n), .Q(
        \l_p_r/counter_r[8] ) );
  NOR2 U246 ( .A(n1137), .B(n208), .Y(n209) );
  MX2 U251 ( .A(n1102), .B(n1103), .S0(n1101), .Y(n214) );
  NOR2B U253 ( .AN(n1103), .B(n1101), .Y(n216) );
  NOR2B U254 ( .AN(n1135), .B(n216), .Y(n217) );
  NOR2 U255 ( .A(n1147), .B(n217), .Y(n218) );
  MX2 U256 ( .A(n211), .B(n1103), .S0(n1136), .Y(n219) );
  NOR2B U257 ( .AN(n1136), .B(n1103), .Y(n220) );
  MX2 U258 ( .A(n211), .B(n1398), .S0(n1137), .Y(n221) );
  MX2 U259 ( .A(n1101), .B(n1137), .S0(n1103), .Y(n222) );
  NOR2 U260 ( .A(n1103), .B(n1101), .Y(n223) );
  MX2 U261 ( .A(n1135), .B(n1134), .S0(n223), .Y(n224) );
  NOR2 U262 ( .A(n1136), .B(n216), .Y(n225) );
  NOR2B U264 ( .AN(n1135), .B(n1163), .Y(n227) );
  NOR2B U265 ( .AN(n211), .B(n1136), .Y(n228) );
  NOR2 U268 ( .A(n1135), .B(n1101), .Y(n231) );
  NOR2B U269 ( .AN(n1103), .B(n1136), .Y(n232) );
  MX2 U270 ( .A(n1100), .B(n1102), .S0(n1135), .Y(n233) );
  MX2 U271 ( .A(n1088), .B(n233), .S0(n1093), .Y(n234) );
  NOR2 U276 ( .A(n211), .B(n217), .Y(n239) );
  MX2 U278 ( .A(n1102), .B(n1392), .S0(n1136), .Y(n241) );
  MX2 U279 ( .A(n1103), .B(n1135), .S0(n1101), .Y(n242) );
  NOR2 U280 ( .A(n1136), .B(n1103), .Y(n243) );
  MX2 U281 ( .A(n1402), .B(n1103), .S0(n1137), .Y(n244) );
  MX2 U282 ( .A(n1137), .B(n1134), .S0(n211), .Y(n245) );
  NOR2B U284 ( .AN(n1136), .B(n223), .Y(n247) );
  NOR2 U285 ( .A(n211), .B(n247), .Y(n248) );
  NOR2B U286 ( .AN(n215), .B(n1089), .Y(n249) );
  MX2 U287 ( .A(n1137), .B(n1134), .S0(n1111), .Y(n250) );
  NOR2B U289 ( .AN(n1135), .B(n1398), .Y(n252) );
  NOR2 U290 ( .A(n223), .B(n252), .Y(n253) );
  NOR2 U291 ( .A(n1392), .B(n217), .Y(n254) );
  NOR2B U292 ( .AN(n236), .B(n211), .Y(n255) );
  MX2 U293 ( .A(n208), .B(n1100), .S0(n1135), .Y(n256) );
  NOR2 U294 ( .A(n212), .B(n1088), .Y(n257) );
  NOR2B U296 ( .AN(n236), .B(n1082), .Y(n259) );
  NOR2B U297 ( .AN(n1140), .B(n1147), .Y(n260) );
  NOR2 U298 ( .A(n1131), .B(n1080), .Y(n261) );
  NOR2 U300 ( .A(n1136), .B(n214), .Y(n263) );
  NOR2 U301 ( .A(n217), .B(n1082), .Y(n264) );
  NOR2B U302 ( .AN(n221), .B(n1132), .Y(n265) );
  NOR2 U304 ( .A(n1133), .B(n1087), .Y(n267) );
  MX2 U305 ( .A(n1137), .B(n1134), .S0(n1103), .Y(n268) );
  MX2 U307 ( .A(n1163), .B(n1101), .S0(n1136), .Y(n270) );
  MX2 U308 ( .A(n1135), .B(n1134), .S0(n1398), .Y(n271) );
  NOR2 U309 ( .A(n209), .B(n220), .Y(n272) );
  NOR2 U310 ( .A(n1131), .B(n1149), .Y(n273) );
  NOR2B U312 ( .AN(n1141), .B(n1411), .Y(n275) );
  NOR2 U313 ( .A(n217), .B(n243), .Y(n276) );
  NOR2B U315 ( .AN(n215), .B(n1088), .Y(n278) );
  MX2 U318 ( .A(n212), .B(n1081), .S0(n1131), .Y(n281) );
  NOR2 U319 ( .A(n1132), .B(n1177), .Y(n282) );
  NOR2 U320 ( .A(n1133), .B(n1077), .Y(n283) );
  NOR2B U321 ( .AN(n261), .B(n247), .Y(n284) );
  NOR2 U322 ( .A(n1131), .B(n1078), .Y(n285) );
  NOR2B U323 ( .AN(n1139), .B(n1149), .Y(n286) );
  MX2 U324 ( .A(n1074), .B(n215), .S0(n1132), .Y(n287) );
  MX2 U326 ( .A(n287), .B(n1396), .S0(\l_p_r/counter_r[2] ), .Y(n289) );
  MX2 U327 ( .A(n288), .B(n258), .S0(n1140), .Y(n290) );
  MX2 U328 ( .A(n285), .B(n283), .S0(n1151), .Y(n291) );
  MX2 U329 ( .A(n289), .B(n290), .S0(n1148), .Y(n292) );
  NOR2 U330 ( .A(n1140), .B(n1149), .Y(n293) );
  AOI222 U331 ( .A0(n1141), .A1(n1411), .B0(n1139), .B1(n1130), .C0(n1150), 
        .C1(n1146), .Y(n294) );
  NOR2B U332 ( .AN(n275), .B(n1090), .Y(n295) );
  MX2 U333 ( .A(n291), .B(n1407), .S0(n1141), .Y(n296) );
  MX2 U334 ( .A(n292), .B(n274), .S0(n1108), .Y(n297) );
  AOI32 U335 ( .A0(n1093), .A1(n1106), .A2(n293), .B0(n1411), .B1(n1108), .Y(
        n298) );
  MX2 U336 ( .A(n294), .B(n295), .S0(n1107), .Y(n299) );
  MX2 U337 ( .A(n267), .B(n296), .S0(n1108), .Y(n300) );
  MX2 U338 ( .A(n297), .B(n298), .S0(n1110), .Y(n301) );
  MX2 U339 ( .A(n299), .B(n300), .S0(n1111), .Y(n302) );
  MX2 U341 ( .A(n1405), .B(n255), .S0(n1133), .Y(n303) );
  AOI32 U342 ( .A0(n1130), .A1(n240), .A2(n1077), .B0(n1132), .B1(n1078), .Y(
        n304) );
  MX2 U343 ( .A(n303), .B(n304), .S0(n1152), .Y(n305) );
  AOI32 U344 ( .A0(n1130), .A1(n230), .A2(n1402), .B0(n1133), .B1(n235), .Y(
        n306) );
  NOR2B U345 ( .AN(n214), .B(n247), .Y(n307) );
  MX2 U346 ( .A(n225), .B(n307), .S0(n1130), .Y(n308) );
  MX2 U347 ( .A(n306), .B(n308), .S0(n1091), .Y(n309) );
  MX2 U348 ( .A(n305), .B(n309), .S0(n1147), .Y(n310) );
  MX2 U349 ( .A(n262), .B(n1089), .S0(n1131), .Y(n311) );
  MX2 U350 ( .A(n248), .B(n1088), .S0(n1132), .Y(n312) );
  MX2 U351 ( .A(n311), .B(n312), .S0(n1151), .Y(n313) );
  NOR2B U352 ( .AN(n258), .B(n1089), .Y(n314) );
  MX2 U353 ( .A(n278), .B(n314), .S0(n1133), .Y(n315) );
  OAI21 U354 ( .A0(\l_p_r/counter_r[2] ), .A1(n315), .B0(n277), .Y(n316) );
  MX2 U355 ( .A(n313), .B(n316), .S0(n1148), .Y(n317) );
  MX2 U356 ( .A(n310), .B(n317), .S0(n1139), .Y(n318) );
  MX2 U357 ( .A(n219), .B(n1404), .S0(n1150), .Y(n319) );
  NOR2B U358 ( .AN(n319), .B(n1131), .Y(n320) );
  NOR2B U359 ( .AN(n1403), .B(n220), .Y(n321) );
  MX2 U360 ( .A(n279), .B(n321), .S0(n1091), .Y(n322) );
  NOR2B U361 ( .AN(n322), .B(n1132), .Y(n323) );
  MX2 U362 ( .A(n320), .B(n323), .S0(n1094), .Y(n324) );
  MX2 U363 ( .A(n252), .B(n1136), .S0(n1090), .Y(n325) );
  MX2 U364 ( .A(n1073), .B(n1403), .S0(n1150), .Y(n326) );
  MX2 U365 ( .A(n325), .B(n326), .S0(n1147), .Y(n327) );
  NOR2B U366 ( .AN(n327), .B(n1133), .Y(n328) );
  MX2 U367 ( .A(n324), .B(n328), .S0(n1140), .Y(n329) );
  MX2 U368 ( .A(n318), .B(n329), .S0(n1107), .Y(n330) );
  NOR2 U369 ( .A(n1140), .B(n1137), .Y(n331) );
  MX2 U371 ( .A(n332), .B(n1411), .S0(n1141), .Y(n333) );
  OAI211 U372 ( .A0(n331), .A1(n333), .B0(n1130), .C0(n1107), .Y(n334) );
  MX2 U373 ( .A(n1100), .B(n1394), .S0(n1152), .Y(n335) );
  MX2 U374 ( .A(n1408), .B(n1178), .S0(n1151), .Y(n336) );
  MX2 U375 ( .A(n335), .B(n336), .S0(n1146), .Y(n337) );
  MX2 U376 ( .A(n1389), .B(n245), .S0(n1091), .Y(n338) );
  MX2 U377 ( .A(n337), .B(n338), .S0(n1139), .Y(n339) );
  MX2 U378 ( .A(n276), .B(n270), .S0(n1152), .Y(n340) );
  NOR2B U379 ( .AN(n1130), .B(n340), .Y(n341) );
  AOI221 U380 ( .A0(n1149), .A1(n280), .B0(n1088), .B1(n280), .C0(n1131), .Y(
        n342) );
  MX2 U381 ( .A(n341), .B(n342), .S0(n1147), .Y(n343) );
  MX2 U383 ( .A(n344), .B(n1400), .S0(n1090), .Y(n345) );
  NOR3 U384 ( .A(n1081), .B(n1132), .C(n1151), .Y(n346) );
  MX2 U385 ( .A(n345), .B(n346), .S0(n1411), .Y(n347) );
  NOR2B U386 ( .AN(n1146), .B(n1130), .Y(n348) );
  NOR2B U387 ( .AN(n347), .B(n348), .Y(n349) );
  MX2 U388 ( .A(n343), .B(n349), .S0(n1140), .Y(n350) );
  OAI2BB2 U389 ( .B0(n334), .B1(n339), .A0N(n1106), .A1N(n350), .Y(n351) );
  MX2 U390 ( .A(n330), .B(n351), .S0(n1110), .Y(\l_p_r/N2850 ) );
  NOR2B U391 ( .AN(n1133), .B(n209), .Y(n352) );
  MX2 U392 ( .A(n1406), .B(n271), .S0(n1131), .Y(n353) );
  MX2 U394 ( .A(n1102), .B(n1075), .S0(n1132), .Y(n355) );
  MX2 U395 ( .A(n1081), .B(n1080), .S0(n1133), .Y(n356) );
  MX2 U396 ( .A(n221), .B(n241), .S0(n1131), .Y(n357) );
  NOR2B U398 ( .AN(n236), .B(n1149), .Y(n359) );
  MX2 U399 ( .A(n263), .B(n211), .S0(n1150), .Y(n360) );
  MX2 U400 ( .A(n223), .B(n1101), .S0(n1137), .Y(n361) );
  NOR2 U402 ( .A(n243), .B(n247), .Y(n363) );
  MX2 U403 ( .A(n353), .B(n354), .S0(n1090), .Y(n364) );
  MX2 U404 ( .A(n355), .B(n274), .S0(\l_p_r/counter_r[2] ), .Y(n365) );
  AOI22 U405 ( .A0(n273), .A1(n1391), .B0(n1149), .B1(n356), .Y(n366) );
  AOI22 U406 ( .A0(n273), .A1(n213), .B0(n1149), .B1(n357), .Y(n367) );
  MX2 U407 ( .A(n276), .B(n1404), .S0(n1151), .Y(n368) );
  MX2 U408 ( .A(n224), .B(n1162), .S0(n1152), .Y(n369) );
  MX2 U409 ( .A(n1102), .B(n1079), .S0(n1091), .Y(n370) );
  NOR2 U410 ( .A(n1131), .B(n1081), .Y(n371) );
  MX2 U411 ( .A(n359), .B(n1149), .S0(n231), .Y(n372) );
  NOR2B U412 ( .AN(n360), .B(n1132), .Y(n373) );
  OAI221 U413 ( .A0(n1152), .A1(n219), .B0(n1149), .B1(n1401), .C0(n1130), .Y(
        n374) );
  MX2 U414 ( .A(n217), .B(n256), .S0(n1151), .Y(n375) );
  MX2 U415 ( .A(n361), .B(n1087), .S0(n1150), .Y(n376) );
  MX2 U416 ( .A(n1161), .B(n363), .S0(n1090), .Y(n377) );
  MX2 U417 ( .A(n364), .B(n365), .S0(n1093), .Y(n378) );
  MX2 U418 ( .A(n366), .B(n367), .S0(n1146), .Y(n379) );
  MX2 U419 ( .A(n1133), .B(n1091), .S0(n275), .Y(n380) );
  MX2 U420 ( .A(n368), .B(n369), .S0(\l_p_r/counter_r[3] ), .Y(n381) );
  MX2 U421 ( .A(n370), .B(n371), .S0(n1146), .Y(n382) );
  AOI32 U422 ( .A0(n372), .A1(n1146), .A2(n1130), .B0(n1411), .B1(n373), .Y(
        n383) );
  MX2 U423 ( .A(n374), .B(n277), .S0(n1094), .Y(n384) );
  MX2 U424 ( .A(n375), .B(n376), .S0(n1093), .Y(n385) );
  MX2 U425 ( .A(n251), .B(n377), .S0(n1148), .Y(n386) );
  MX2 U426 ( .A(n378), .B(n379), .S0(n1141), .Y(n387) );
  NOR2B U427 ( .AN(n1108), .B(n380), .Y(n388) );
  MX2 U428 ( .A(n381), .B(n382), .S0(n1139), .Y(n389) );
  MX2 U429 ( .A(n383), .B(n384), .S0(n1140), .Y(n390) );
  MX2 U430 ( .A(n385), .B(n386), .S0(n1141), .Y(n391) );
  AOI211 U431 ( .A0(n1151), .A1(n260), .B0(n1131), .C0(n1107), .Y(n392) );
  OAI2BB2 U432 ( .B0(n1107), .B1(n387), .A0N(n388), .A1N(n389), .Y(n393) );
  OAI2BB2 U433 ( .B0(n390), .B1(n1106), .A0N(n391), .A1N(n392), .Y(n394) );
  MX2 U434 ( .A(n393), .B(n394), .S0(n1111), .Y(\l_p_r/N2851 ) );
  MX2 U435 ( .A(n1100), .B(n1398), .S0(n1132), .Y(n395) );
  MX2 U436 ( .A(n1135), .B(n1134), .S0(n1133), .Y(n396) );
  MX2 U437 ( .A(n214), .B(n1392), .S0(n1135), .Y(n397) );
  MX2 U438 ( .A(n395), .B(n211), .S0(n396), .Y(n398) );
  NOR2B U439 ( .AN(n261), .B(n213), .Y(n399) );
  MX2 U440 ( .A(n262), .B(n1080), .S0(n1131), .Y(n400) );
  MX2 U441 ( .A(n263), .B(n1089), .S0(n1132), .Y(n401) );
  MX2 U442 ( .A(n264), .B(n243), .S0(n1133), .Y(n402) );
  MX2 U443 ( .A(n1163), .B(n266), .S0(n1131), .Y(n403) );
  NOR2B U444 ( .AN(n213), .B(n1132), .Y(n404) );
  MX2 U445 ( .A(n1088), .B(n1404), .S0(n1090), .Y(n405) );
  MX2 U446 ( .A(n239), .B(n270), .S0(n1150), .Y(n406) );
  MX2 U447 ( .A(n254), .B(n259), .S0(n1152), .Y(n407) );
  MX2 U448 ( .A(n271), .B(n1136), .S0(n1151), .Y(n408) );
  MX2 U449 ( .A(n272), .B(n1087), .S0(n1091), .Y(n409) );
  MX2 U450 ( .A(n1405), .B(n211), .S0(n1152), .Y(n410) );
  MX2 U451 ( .A(n1088), .B(n397), .S0(n1091), .Y(n411) );
  MX2 U452 ( .A(n1103), .B(n213), .S0(n1150), .Y(n412) );
  MX2 U453 ( .A(n398), .B(n399), .S0(n1090), .Y(n413) );
  MX2 U454 ( .A(n400), .B(n401), .S0(\l_p_r/counter_r[2] ), .Y(n414) );
  MX2 U455 ( .A(n402), .B(n265), .S0(n1151), .Y(n415) );
  MX2 U456 ( .A(n403), .B(n404), .S0(n1152), .Y(n416) );
  NOR2B U457 ( .AN(n230), .B(n1133), .Y(n417) );
  NOR2B U458 ( .AN(n405), .B(n1131), .Y(n418) );
  MX2 U459 ( .A(n406), .B(n407), .S0(n1094), .Y(n419) );
  MX2 U460 ( .A(n408), .B(n409), .S0(n1093), .Y(n420) );
  NOR2B U461 ( .AN(n410), .B(n1132), .Y(n421) );
  NOR2B U462 ( .AN(n411), .B(n1133), .Y(n422) );
  AOI32 U463 ( .A0(n220), .A1(n1147), .A2(n273), .B0(n412), .B1(n1411), .Y(
        n423) );
  NOR2B U464 ( .AN(n1131), .B(n1094), .Y(n424) );
  MX2 U465 ( .A(n413), .B(n414), .S0(n1148), .Y(n425) );
  MX2 U466 ( .A(n415), .B(n416), .S0(n1147), .Y(n426) );
  AOI32 U467 ( .A0(n417), .A1(n1093), .A2(n237), .B0(n1411), .B1(n418), .Y(
        n427) );
  AOI32 U468 ( .A0(n267), .A1(n1141), .A2(n1411), .B0(n1149), .B1(n1139), .Y(
        n428) );
  MX2 U469 ( .A(n269), .B(n1395), .S0(n1148), .Y(n429) );
  MX2 U470 ( .A(n419), .B(n420), .S0(n1139), .Y(n430) );
  MX2 U471 ( .A(n421), .B(n422), .S0(n1094), .Y(n431) );
  NOR2 U472 ( .A(n423), .B(n424), .Y(n432) );
  MX2 U473 ( .A(n425), .B(n426), .S0(n1140), .Y(n433) );
  OAI22 U474 ( .A0(n1140), .A1(n427), .B0(n428), .B1(n429), .Y(n434) );
  NOR2 U475 ( .A(n1132), .B(n430), .Y(n435) );
  MX2 U476 ( .A(n431), .B(n432), .S0(n1141), .Y(n436) );
  MX2 U477 ( .A(n433), .B(n434), .S0(n1108), .Y(n437) );
  MX2 U478 ( .A(n435), .B(n436), .S0(n1107), .Y(n438) );
  MX2 U479 ( .A(n437), .B(n438), .S0(n1110), .Y(\l_p_r/N2852 ) );
  NOR2B U480 ( .AN(n1074), .B(n213), .Y(n439) );
  MX2 U481 ( .A(n1134), .B(n1137), .S0(n1101), .Y(n440) );
  NOR2B U482 ( .AN(n1110), .B(n1398), .Y(n441) );
  MX2 U483 ( .A(n1176), .B(n208), .S0(n1111), .Y(n442) );
  MX2 U484 ( .A(n439), .B(n248), .S0(n1110), .Y(n443) );
  MX2 U485 ( .A(n212), .B(n1089), .S0(n1111), .Y(n444) );
  MX2 U486 ( .A(n440), .B(n249), .S0(n1110), .Y(n445) );
  MX2 U487 ( .A(n1176), .B(n441), .S0(n250), .Y(n446) );
  MX2 U488 ( .A(n1102), .B(n442), .S0(n250), .Y(n447) );
  AOI211 U489 ( .A0(n1111), .A1(n1404), .B0(n1079), .C0(n1084), .Y(n448) );
  MX2 U490 ( .A(n1176), .B(n1078), .S0(n1111), .Y(n449) );
  MX2 U491 ( .A(n1387), .B(n251), .S0(n1110), .Y(n450) );
  MX2 U492 ( .A(n253), .B(n244), .S0(n1111), .Y(n451) );
  MX2 U493 ( .A(n235), .B(n254), .S0(n1110), .Y(n452) );
  MX2 U494 ( .A(n255), .B(n256), .S0(n1111), .Y(n453) );
  MX2 U495 ( .A(n1397), .B(n257), .S0(n1110), .Y(n454) );
  AOI211 U496 ( .A0(n1110), .A1(n258), .B0(n1081), .C0(n1084), .Y(n455) );
  MX2 U497 ( .A(n1177), .B(n1389), .S0(n1111), .Y(n456) );
  MX2 U498 ( .A(n1134), .B(n243), .S0(n1110), .Y(n457) );
  MX2 U500 ( .A(n443), .B(n444), .S0(n1108), .Y(n459) );
  MX2 U501 ( .A(n445), .B(n446), .S0(n1107), .Y(n460) );
  MX2 U502 ( .A(n447), .B(n448), .S0(n1108), .Y(n461) );
  MX2 U503 ( .A(n449), .B(n450), .S0(n1107), .Y(n462) );
  MX2 U504 ( .A(n451), .B(n452), .S0(n1108), .Y(n463) );
  MX2 U505 ( .A(n453), .B(n454), .S0(n1107), .Y(n464) );
  MX2 U506 ( .A(n455), .B(n456), .S0(n1108), .Y(n465) );
  MX2 U507 ( .A(n457), .B(n458), .S0(n1107), .Y(n466) );
  MX2 U508 ( .A(n459), .B(n460), .S0(n1139), .Y(n467) );
  MX2 U509 ( .A(n461), .B(n462), .S0(n1140), .Y(n468) );
  MX2 U510 ( .A(n463), .B(n464), .S0(n1141), .Y(n469) );
  MX2 U511 ( .A(n465), .B(n466), .S0(n1139), .Y(n470) );
  MX2 U512 ( .A(n1391), .B(n1089), .S0(n1140), .Y(n471) );
  MX2 U513 ( .A(n1080), .B(n259), .S0(n1141), .Y(n472) );
  MX2 U514 ( .A(n467), .B(n468), .S0(n1091), .Y(n473) );
  MX2 U515 ( .A(n469), .B(n470), .S0(n1151), .Y(n474) );
  MX2 U516 ( .A(n471), .B(n1082), .S0(n1150), .Y(n475) );
  MX2 U517 ( .A(n472), .B(n1089), .S0(n1091), .Y(n476) );
  MX2 U519 ( .A(n473), .B(n474), .S0(n1147), .Y(n478) );
  MX2 U520 ( .A(n475), .B(n476), .S0(n1146), .Y(n479) );
  AOI211 U521 ( .A0(n1150), .A1(n260), .B0(n1111), .C0(n477), .Y(n480) );
  OAI2BB2 U522 ( .B0(n1133), .B1(n478), .A0N(n479), .A1N(n480), .Y(
        \l_p_r/N2853 ) );
  MX2 U523 ( .A(n1101), .B(n1398), .S0(n1136), .Y(n481) );
  MX2 U524 ( .A(n481), .B(n1135), .S0(n1411), .Y(n482) );
  NOR2B U525 ( .AN(n1149), .B(n482), .Y(n483) );
  MX2 U526 ( .A(n1077), .B(n284), .S0(n1090), .Y(n484) );
  NOR2B U527 ( .AN(n484), .B(n1141), .Y(n485) );
  MX2 U528 ( .A(n1102), .B(n1399), .S0(n1132), .Y(n486) );
  MX2 U529 ( .A(n1134), .B(n1080), .S0(n1133), .Y(n487) );
  MX2 U530 ( .A(n486), .B(n487), .S0(n1147), .Y(n488) );
  MX2 U531 ( .A(n1393), .B(n1089), .S0(n1131), .Y(n489) );
  MX2 U532 ( .A(n281), .B(n489), .S0(n1093), .Y(n490) );
  MX2 U533 ( .A(n488), .B(n490), .S0(n1150), .Y(n491) );
  MX2 U534 ( .A(n1082), .B(n1408), .S0(n1132), .Y(n492) );
  OAI2BB2 U535 ( .B0(n492), .B1(n1411), .A0N(n259), .A1N(n1130), .Y(n493) );
  MX2 U536 ( .A(n1163), .B(n216), .S0(n1411), .Y(n494) );
  MX2 U537 ( .A(n1411), .B(n1093), .S0(n1137), .Y(n495) );
  MX2 U538 ( .A(n494), .B(n1402), .S0(n495), .Y(n496) );
  MX2 U539 ( .A(n1077), .B(n258), .S0(n1146), .Y(n497) );
  NOR2B U540 ( .AN(n497), .B(n1130), .Y(n498) );
  NOR2B U541 ( .AN(n496), .B(n498), .Y(n499) );
  MX2 U542 ( .A(n493), .B(n499), .S0(n1149), .Y(n500) );
  MX2 U543 ( .A(n491), .B(n500), .S0(n1139), .Y(n501) );
  MX2 U544 ( .A(n259), .B(n1136), .S0(\l_p_r/counter_r[3] ), .Y(n502) );
  MX2 U545 ( .A(n1082), .B(n502), .S0(n1152), .Y(n503) );
  MX2 U546 ( .A(n1080), .B(n1406), .S0(n1146), .Y(n504) );
  AOI21 U547 ( .A0(n504), .A1(n1090), .B0(n483), .Y(n505) );
  MX2 U548 ( .A(n503), .B(n505), .S0(n1140), .Y(n506) );
  NOR2B U549 ( .AN(n506), .B(n1131), .Y(n507) );
  MX2 U550 ( .A(n501), .B(n507), .S0(n1108), .Y(n508) );
  AOI32 U551 ( .A0(n1130), .A1(n272), .A2(n1146), .B0(n1388), .B1(n1130), .Y(
        n509) );
  MX2 U552 ( .A(n280), .B(n1390), .S0(n1094), .Y(n510) );
  OAI2BB2 U553 ( .B0(n1090), .B1(n509), .A0N(n273), .A1N(n510), .Y(n511) );
  AOI32 U555 ( .A0(n485), .A1(n1130), .A2(n1084), .B0(n512), .B1(n485), .Y(
        n513) );
  AOI221 U556 ( .A0(n1411), .A1(n1130), .B0(n1401), .B1(n1130), .C0(n1150), 
        .Y(n514) );
  AOI2BB2 U557 ( .B0(n1139), .B1(n511), .A0N(n513), .A1N(n514), .Y(n515) );
  MX2 U558 ( .A(n248), .B(n244), .S0(n1094), .Y(n516) );
  NOR2B U559 ( .AN(n1406), .B(n213), .Y(n517) );
  MX2 U560 ( .A(n257), .B(n517), .S0(n1148), .Y(n518) );
  MX2 U561 ( .A(n516), .B(n518), .S0(n1151), .Y(n519) );
  MX2 U562 ( .A(n249), .B(n1389), .S0(n1093), .Y(n520) );
  MX2 U563 ( .A(n520), .B(n269), .S0(n1091), .Y(n521) );
  MX2 U564 ( .A(n519), .B(n521), .S0(n1141), .Y(n522) );
  OAI221 U565 ( .A0(n1410), .A1(n1093), .B0(n286), .B1(n1130), .C0(n1106), .Y(
        n523) );
  OAI22 U566 ( .A0(n515), .A1(n1106), .B0(n522), .B1(n523), .Y(n524) );
  MX2 U567 ( .A(n508), .B(n524), .S0(n1111), .Y(\l_p_r/N2854 ) );
  MX2 U568 ( .A(n1101), .B(n214), .S0(n1135), .Y(n525) );
  AOI32 U569 ( .A0(n1077), .A1(n1132), .A2(n258), .B0(n1103), .B1(n1130), .Y(
        n526) );
  NOR2 U570 ( .A(n1133), .B(n237), .Y(n527) );
  MX2 U571 ( .A(n251), .B(n1137), .S0(n1133), .Y(n528) );
  MX2 U572 ( .A(n233), .B(n1163), .S0(n1131), .Y(n529) );
  MX2 U573 ( .A(n268), .B(n258), .S0(n1132), .Y(n530) );
  MX2 U574 ( .A(n266), .B(n1135), .S0(n1093), .Y(n531) );
  MX2 U575 ( .A(n235), .B(n525), .S0(n1148), .Y(n532) );
  AOI32 U576 ( .A0(n1073), .A1(n1411), .A2(n280), .B0(n1148), .B1(n241), .Y(
        n533) );
  NOR2 U577 ( .A(n1079), .B(n1084), .Y(n534) );
  MX2 U578 ( .A(n526), .B(n527), .S0(n1147), .Y(n535) );
  MX2 U579 ( .A(n281), .B(n528), .S0(n1148), .Y(n536) );
  MX2 U580 ( .A(n529), .B(n530), .S0(n1094), .Y(n537) );
  AOI32 U581 ( .A0(n1148), .A1(n1151), .A2(n1081), .B0(n1130), .B1(n1150), .Y(
        n538) );
  MX2 U582 ( .A(n255), .B(n224), .S0(n1147), .Y(n539) );
  MX2 U583 ( .A(n282), .B(n283), .S0(n1146), .Y(n540) );
  NOR2B U584 ( .AN(n531), .B(n1131), .Y(n541) );
  MX2 U585 ( .A(n1388), .B(n1077), .S0(n1147), .Y(n542) );
  MX2 U586 ( .A(n284), .B(n285), .S0(n1093), .Y(n543) );
  MX2 U587 ( .A(n1102), .B(n1148), .S0(n1101), .Y(n544) );
  OAI211 U588 ( .A0(n1094), .A1(n236), .B0(n1130), .C0(n1149), .Y(n545) );
  MX2 U589 ( .A(n532), .B(n533), .S0(n1152), .Y(n546) );
  AOI32 U590 ( .A0(n1178), .A1(n1147), .A2(n1406), .B0(n534), .B1(n1411), .Y(
        n547) );
  MX2 U591 ( .A(n254), .B(n241), .S0(n1146), .Y(n548) );
  MX2 U592 ( .A(n1082), .B(n1088), .S0(\l_p_r/counter_r[3] ), .Y(n549) );
  NOR2 U593 ( .A(n1140), .B(n1091), .Y(n550) );
  MX2 U594 ( .A(n535), .B(n536), .S0(n1090), .Y(n551) );
  OAI22 U595 ( .A0(n1152), .A1(n537), .B0(n538), .B1(n539), .Y(n552) );
  MX2 U596 ( .A(n540), .B(n541), .S0(n1150), .Y(n553) );
  AOI211 U597 ( .A0(n1152), .A1(n542), .B0(n1132), .C0(n483), .Y(n554) );
  AOI2BB2 U598 ( .B0(n1152), .B1(n543), .A0N(n544), .A1N(n545), .Y(n555) );
  MX2 U600 ( .A(n282), .B(n547), .S0(n1090), .Y(n557) );
  MX2 U601 ( .A(n548), .B(n549), .S0(\l_p_r/counter_r[2] ), .Y(n558) );
  MX2 U602 ( .A(n1133), .B(n1147), .S0(n550), .Y(n559) );
  MX2 U603 ( .A(n551), .B(n552), .S0(n1139), .Y(n560) );
  MX2 U604 ( .A(n553), .B(n554), .S0(n1140), .Y(n561) );
  MX2 U605 ( .A(n555), .B(n556), .S0(n1141), .Y(n562) );
  MX2 U606 ( .A(n557), .B(n558), .S0(n1139), .Y(n563) );
  NOR2B U607 ( .AN(n1106), .B(n559), .Y(n564) );
  MX2 U608 ( .A(n560), .B(n561), .S0(n1107), .Y(n565) );
  OAI2BB2 U609 ( .B0(n562), .B1(n1106), .A0N(n563), .A1N(n564), .Y(n566) );
  MX2 U610 ( .A(n565), .B(n566), .S0(n1110), .Y(\l_p_r/N2855 ) );
  NOR2B U611 ( .AN(n215), .B(n216), .Y(n567) );
  MX2 U612 ( .A(n1081), .B(n1084), .S0(n1146), .Y(n568) );
  NOR2B U613 ( .AN(n1148), .B(n217), .Y(n569) );
  MX2 U614 ( .A(n239), .B(n1405), .S0(n1094), .Y(n570) );
  OAI31 U615 ( .A0(n1079), .A1(n1084), .A2(n1411), .B0(n240), .Y(n571) );
  MX2 U616 ( .A(n241), .B(n220), .S0(n1094), .Y(n572) );
  MX2 U617 ( .A(n221), .B(n242), .S0(n1148), .Y(n573) );
  MX2 U618 ( .A(n224), .B(n243), .S0(n1094), .Y(n574) );
  MX2 U619 ( .A(n219), .B(n215), .S0(n1093), .Y(n575) );
  MX2 U621 ( .A(n230), .B(n1087), .S0(n1148), .Y(n577) );
  MX2 U622 ( .A(n1403), .B(n245), .S0(n1147), .Y(n578) );
  MX2 U623 ( .A(n1136), .B(n1080), .S0(n1148), .Y(n579) );
  OAI2BB1 U624 ( .A0N(n1093), .A1N(n236), .B0(n1077), .Y(n580) );
  MX2 U625 ( .A(n222), .B(n1134), .S0(n1094), .Y(n581) );
  AOI32 U626 ( .A0(n214), .A1(n1411), .A2(n230), .B0(n239), .B1(n1146), .Y(
        n582) );
  MX2 U627 ( .A(n1411), .B(n1146), .S0(n1079), .Y(n583) );
  MX2 U628 ( .A(n244), .B(n567), .S0(n1411), .Y(n584) );
  MX2 U629 ( .A(n568), .B(n569), .S0(n1151), .Y(n585) );
  MX2 U630 ( .A(n570), .B(n571), .S0(n1152), .Y(n586) );
  MX2 U631 ( .A(n218), .B(n572), .S0(n1091), .Y(n587) );
  MX2 U632 ( .A(n573), .B(n574), .S0(n1151), .Y(n588) );
  OAI32 U633 ( .A0(n1090), .A1(n1147), .A2(n239), .B0(n575), .B1(n1149), .Y(
        n589) );
  MX2 U634 ( .A(n576), .B(n577), .S0(n1150), .Y(n590) );
  MX2 U635 ( .A(n578), .B(n579), .S0(\l_p_r/counter_r[2] ), .Y(n591) );
  MX2 U636 ( .A(n580), .B(n581), .S0(n1090), .Y(n592) );
  MX2 U637 ( .A(n582), .B(n583), .S0(n1150), .Y(n593) );
  MX2 U638 ( .A(n234), .B(n584), .S0(n1152), .Y(n594) );
  MX2 U639 ( .A(n585), .B(n586), .S0(n1140), .Y(n595) );
  MX2 U640 ( .A(n587), .B(n588), .S0(n1141), .Y(n596) );
  MX2 U641 ( .A(n589), .B(n590), .S0(n1139), .Y(n597) );
  MX2 U642 ( .A(n591), .B(n592), .S0(n1140), .Y(n598) );
  MX2 U643 ( .A(n593), .B(n594), .S0(n1141), .Y(n599) );
  MX2 U644 ( .A(n595), .B(n596), .S0(n1108), .Y(n600) );
  NOR2 U645 ( .A(n1108), .B(n597), .Y(n601) );
  MX2 U646 ( .A(n598), .B(n599), .S0(n1107), .Y(n602) );
  MX2 U647 ( .A(n600), .B(n601), .S0(n1133), .Y(n603) );
  NOR2B U648 ( .AN(n602), .B(n1131), .Y(n604) );
  MX2 U649 ( .A(n603), .B(n604), .S0(n1111), .Y(\l_p_r/N2856 ) );
  MX2 U650 ( .A(n1398), .B(n1402), .S0(n1136), .Y(n605) );
  MX2 U651 ( .A(n1103), .B(n1176), .S0(n1137), .Y(n606) );
  NOR2B U652 ( .AN(n236), .B(n216), .Y(n607) );
  MX2 U653 ( .A(n1402), .B(n1398), .S0(n1135), .Y(n608) );
  NOR2B U654 ( .AN(n209), .B(n1094), .Y(n609) );
  MX2 U655 ( .A(n212), .B(n213), .S0(n1147), .Y(n610) );
  OAI222 U656 ( .A0(n1137), .A1(n1103), .B0(n1135), .B1(n1094), .C0(n215), 
        .C1(n1411), .Y(n611) );
  AOI211 U657 ( .A0(n1136), .A1(n1101), .B0(n1094), .C0(n1103), .Y(n612) );
  MX2 U658 ( .A(n219), .B(n220), .S0(n1146), .Y(n613) );
  MX2 U659 ( .A(n221), .B(n222), .S0(n1147), .Y(n614) );
  MX2 U660 ( .A(n224), .B(n225), .S0(n1093), .Y(n615) );
  MX2 U661 ( .A(n605), .B(n1089), .S0(n1146), .Y(n616) );
  NOR2B U662 ( .AN(n606), .B(n1146), .Y(n617) );
  MX2 U663 ( .A(n1082), .B(n1084), .S0(\l_p_r/counter_r[3] ), .Y(n618) );
  MX2 U664 ( .A(n213), .B(n1079), .S0(n1146), .Y(n619) );
  MX2 U665 ( .A(n235), .B(n1074), .S0(n1094), .Y(n620) );
  MX2 U666 ( .A(n1137), .B(n1403), .S0(\l_p_r/counter_r[3] ), .Y(n621) );
  MX2 U667 ( .A(n237), .B(n607), .S0(n1148), .Y(n622) );
  MX2 U668 ( .A(n1087), .B(n1134), .S0(n1093), .Y(n623) );
  MX2 U669 ( .A(n1077), .B(n230), .S0(n1093), .Y(n624) );
  MX2 U670 ( .A(n1411), .B(n1093), .S0(n231), .Y(n625) );
  MX2 U671 ( .A(n608), .B(n1387), .S0(n1148), .Y(n626) );
  MX2 U672 ( .A(n609), .B(n610), .S0(n1151), .Y(n627) );
  MX2 U673 ( .A(n611), .B(n218), .S0(n1091), .Y(n628) );
  MX2 U674 ( .A(n612), .B(n613), .S0(n1152), .Y(n629) );
  MX2 U675 ( .A(n614), .B(n615), .S0(n1091), .Y(n630) );
  MX2 U676 ( .A(n616), .B(n617), .S0(n1150), .Y(n631) );
  MX2 U677 ( .A(n618), .B(n619), .S0(n1090), .Y(n632) );
  MX2 U678 ( .A(n620), .B(n621), .S0(\l_p_r/counter_r[2] ), .Y(n633) );
  MX2 U679 ( .A(n622), .B(n623), .S0(n1151), .Y(n634) );
  MX2 U680 ( .A(n624), .B(n625), .S0(n1152), .Y(n635) );
  MX2 U681 ( .A(n234), .B(n626), .S0(n1091), .Y(n636) );
  MX2 U682 ( .A(n627), .B(n628), .S0(n1139), .Y(n637) );
  MX2 U683 ( .A(n629), .B(n630), .S0(n1140), .Y(n638) );
  MX2 U684 ( .A(n631), .B(n632), .S0(n1141), .Y(n639) );
  MX2 U685 ( .A(n633), .B(n634), .S0(n1139), .Y(n640) );
  MX2 U686 ( .A(n635), .B(n636), .S0(n1140), .Y(n641) );
  MX2 U687 ( .A(n637), .B(n638), .S0(n1108), .Y(n642) );
  NOR2B U688 ( .AN(n639), .B(n1107), .Y(n643) );
  MX2 U689 ( .A(n640), .B(n641), .S0(n1107), .Y(n644) );
  MX2 U690 ( .A(n642), .B(n643), .S0(n1131), .Y(n645) );
  NOR2B U691 ( .AN(n644), .B(n1132), .Y(n646) );
  MX2 U692 ( .A(n645), .B(n646), .S0(n1110), .Y(\l_p_r/N2857 ) );
  MX2 U695 ( .A(n1155), .B(n1153), .S0(n1143), .Y(n649) );
  NOR2B U700 ( .AN(n1105), .B(n1086), .Y(n654) );
  MX2 U701 ( .A(n1099), .B(n1105), .S0(n1120), .Y(n655) );
  NOR2B U702 ( .AN(n1120), .B(n1099), .Y(n656) );
  MX2 U703 ( .A(n1105), .B(n1104), .S0(n1086), .Y(n657) );
  NOR2 U705 ( .A(n1097), .B(n658), .Y(n659) );
  MX2 U706 ( .A(n1105), .B(n1099), .S0(n1121), .Y(n660) );
  MX2 U707 ( .A(n660), .B(n1099), .S0(\r_p_r/counter_r[4] ), .Y(n661) );
  NOR2 U709 ( .A(n1121), .B(n662), .Y(n663) );
  MX2 U711 ( .A(n1105), .B(n1385), .S0(n1119), .Y(n665) );
  MX2 U713 ( .A(n1105), .B(n1158), .S0(n1120), .Y(n667) );
  MX2 U715 ( .A(n1104), .B(n1386), .S0(n1121), .Y(n669) );
  NOR2B U716 ( .AN(n1119), .B(n1382), .Y(n670) );
  NOR2 U717 ( .A(n1097), .B(n667), .Y(n671) );
  MX2 U719 ( .A(n1092), .B(n1099), .S0(n1096), .Y(n673) );
  MX2 U720 ( .A(n651), .B(n1105), .S0(n1119), .Y(n674) );
  MX2 U721 ( .A(n1383), .B(n1104), .S0(n1120), .Y(n675) );
  MX2 U723 ( .A(n1372), .B(n676), .S0(n1097), .Y(n677) );
  MX2 U724 ( .A(n1120), .B(n1086), .S0(n1105), .Y(n678) );
  MX2 U725 ( .A(n678), .B(n1104), .S0(n1095), .Y(n679) );
  NOR2 U726 ( .A(n1121), .B(n1105), .Y(n680) );
  MX2 U728 ( .A(n1386), .B(n1385), .S0(n1121), .Y(n682) );
  NOR2B U729 ( .AN(n1119), .B(n662), .Y(n683) );
  NOR2B U730 ( .AN(n1120), .B(n1158), .Y(n684) );
  NOR2B U733 ( .AN(n1121), .B(n1386), .Y(n687) );
  MX2 U735 ( .A(n1374), .B(n688), .S0(n1097), .Y(n689) );
  MX2 U736 ( .A(n1105), .B(n1086), .S0(n1119), .Y(n690) );
  MX2 U738 ( .A(n1158), .B(n1086), .S0(n1120), .Y(n692) );
  MX2 U741 ( .A(n1383), .B(n651), .S0(n1121), .Y(n697) );
  OAI221 U742 ( .A0(n1095), .A1(n697), .B0(n1142), .B1(n1119), .C0(n1153), .Y(
        n698) );
  MX2 U744 ( .A(n1386), .B(n1158), .S0(n1143), .Y(n700) );
  NOR2B U745 ( .AN(n1120), .B(n651), .Y(n701) );
  MX2 U746 ( .A(n701), .B(n1366), .S0(n1096), .Y(n702) );
  NOR2B U747 ( .AN(n686), .B(n1386), .Y(n703) );
  NOR2 U748 ( .A(n703), .B(n1142), .Y(n704) );
  NOR2 U749 ( .A(n1144), .B(n1158), .Y(n705) );
  MX2 U750 ( .A(n1382), .B(n1085), .S0(n1119), .Y(n706) );
  NOR2B U751 ( .AN(n1105), .B(n1121), .Y(n707) );
  NOR2B U752 ( .AN(n1119), .B(n1098), .Y(n708) );
  NOR2B U753 ( .AN(n663), .B(n1096), .Y(n709) );
  MX2 U754 ( .A(n665), .B(n685), .S0(n1097), .Y(n710) );
  MX2 U755 ( .A(n1144), .B(n1142), .S0(n1120), .Y(n711) );
  NOR2 U756 ( .A(\r_p_r/counter_r[4] ), .B(n674), .Y(n712) );
  NOR2 U757 ( .A(n657), .B(n684), .Y(n713) );
  NOR2 U758 ( .A(n1143), .B(n1379), .Y(n714) );
  NOR2 U763 ( .A(n1120), .B(n1099), .Y(n719) );
  NOR2 U764 ( .A(n1121), .B(n657), .Y(n720) );
  MX2 U765 ( .A(n701), .B(n720), .S0(n1144), .Y(n721) );
  NOR2 U766 ( .A(n680), .B(n701), .Y(n722) );
  OAI21 U770 ( .A0(n1113), .A1(n1379), .B0(n1116), .Y(n726) );
  MX2 U771 ( .A(n663), .B(n715), .S0(n1124), .Y(n727) );
  MX2 U772 ( .A(n701), .B(n1375), .S0(n1123), .Y(n728) );
  MX2 U774 ( .A(n1156), .B(n1153), .S0(n1124), .Y(n730) );
  MX2 U775 ( .A(n1382), .B(n727), .S0(n1154), .Y(n731) );
  MX2 U776 ( .A(n1092), .B(n728), .S0(n1157), .Y(n732) );
  MX2 U777 ( .A(n708), .B(n683), .S0(n1127), .Y(n733) );
  MX2 U778 ( .A(n1129), .B(n1125), .S0(n1156), .Y(n734) );
  AOI33 U779 ( .A0(n1156), .A1(n1123), .A2(n715), .B0(n1092), .B1(n1122), .B2(
        n1153), .Y(n735) );
  MX2 U780 ( .A(n1117), .B(n729), .S0(n730), .Y(n736) );
  AOI33 U781 ( .A0(n1116), .A1(n1124), .A2(n1153), .B0(n1156), .B1(n1122), 
        .B2(n1115), .Y(n737) );
  NOR2 U782 ( .A(n1117), .B(n1154), .Y(n738) );
  MX2 U783 ( .A(n731), .B(n732), .S0(n1128), .Y(n739) );
  MX2 U784 ( .A(n733), .B(n1380), .S0(n734), .Y(n740) );
  MX2 U785 ( .A(n715), .B(n1386), .S0(n1123), .Y(n741) );
  NOR2 U786 ( .A(n735), .B(n1116), .Y(n742) );
  MX2 U787 ( .A(n736), .B(n737), .S0(n1144), .Y(n743) );
  AOI32 U788 ( .A0(n1126), .A1(n1142), .A2(n738), .B0(n1125), .B1(n1097), .Y(
        n744) );
  MX2 U789 ( .A(n739), .B(n740), .S0(n1097), .Y(n745) );
  MX2 U790 ( .A(n741), .B(n742), .S0(n1097), .Y(n746) );
  MX2 U791 ( .A(n743), .B(n744), .S0(n1113), .Y(n747) );
  MX2 U792 ( .A(n745), .B(n746), .S0(n1114), .Y(n748) );
  MX2 U794 ( .A(n657), .B(n1105), .S0(n1121), .Y(n749) );
  NOR2 U795 ( .A(n1092), .B(n715), .Y(n750) );
  MX2 U796 ( .A(n1105), .B(n1099), .S0(n1113), .Y(n751) );
  MX2 U797 ( .A(n1119), .B(n1118), .S0(n1114), .Y(n752) );
  NOR2B U798 ( .AN(n693), .B(n715), .Y(n753) );
  MX2 U799 ( .A(n1105), .B(n1383), .S0(n1113), .Y(n754) );
  NOR2B U800 ( .AN(n697), .B(n1114), .Y(n755) );
  MX2 U801 ( .A(n680), .B(n1379), .S0(n1114), .Y(n756) );
  MX2 U802 ( .A(n658), .B(n674), .S0(n1113), .Y(n757) );
  MX2 U803 ( .A(n749), .B(n1370), .S0(n1114), .Y(n758) );
  MX2 U804 ( .A(n666), .B(n750), .S0(n1113), .Y(n759) );
  MX2 U806 ( .A(n751), .B(n1158), .S0(n752), .Y(n761) );
  NOR2B U807 ( .AN(n688), .B(n1113), .Y(n762) );
  MX2 U808 ( .A(n713), .B(n1381), .S0(n1114), .Y(n763) );
  MX2 U809 ( .A(n703), .B(n1180), .S0(n1113), .Y(n764) );
  MX2 U811 ( .A(n1382), .B(n720), .S0(n1114), .Y(n766) );
  NOR2B U812 ( .AN(n713), .B(n1114), .Y(n767) );
  MX2 U813 ( .A(n1104), .B(n670), .S0(n1113), .Y(n768) );
  NOR2 U814 ( .A(n1113), .B(n651), .Y(n769) );
  MX2 U815 ( .A(n715), .B(n753), .S0(n1117), .Y(n770) );
  MX2 U816 ( .A(n665), .B(n1386), .S0(n1116), .Y(n771) );
  MX2 U817 ( .A(n754), .B(n755), .S0(n1117), .Y(n772) );
  OAI32 U818 ( .A0(n1115), .A1(n1114), .A2(n707), .B0(n1117), .B1(n756), .Y(
        n773) );
  MX2 U819 ( .A(n757), .B(n725), .S0(n1116), .Y(n774) );
  MX2 U820 ( .A(n1158), .B(n1385), .S0(n1117), .Y(n775) );
  NOR2 U821 ( .A(n1113), .B(n1369), .Y(n776) );
  AOI21 U822 ( .A0(n1116), .A1(n670), .B0(n1114), .Y(n777) );
  MX2 U823 ( .A(n758), .B(n725), .S0(n1116), .Y(n778) );
  MX2 U824 ( .A(n759), .B(n760), .S0(n1117), .Y(n779) );
  MX2 U825 ( .A(n761), .B(n762), .S0(n1116), .Y(n780) );
  NOR2B U826 ( .AN(n726), .B(n763), .Y(n781) );
  MX2 U827 ( .A(n764), .B(n765), .S0(n1117), .Y(n782) );
  MX2 U828 ( .A(n766), .B(n767), .S0(n1116), .Y(n783) );
  MX2 U829 ( .A(n768), .B(n769), .S0(n1117), .Y(n784) );
  NOR2B U830 ( .AN(n770), .B(n1113), .Y(n785) );
  NOR2B U831 ( .AN(n771), .B(n1114), .Y(n786) );
  MX2 U832 ( .A(n772), .B(n773), .S0(n1157), .Y(n787) );
  OAI32 U833 ( .A0(n1153), .A1(n724), .A2(n1085), .B0(n1155), .B1(n774), .Y(
        n788) );
  NOR2B U834 ( .AN(n1155), .B(n775), .Y(n789) );
  AOI32 U835 ( .A0(n776), .A1(n1153), .A2(n726), .B0(n1155), .B1(n777), .Y(
        n790) );
  MX2 U836 ( .A(n778), .B(n779), .S0(\r_p_r/counter_r[5] ), .Y(n791) );
  MX2 U837 ( .A(n780), .B(n781), .S0(n1156), .Y(n792) );
  OAI32 U838 ( .A0(n1157), .A1(n1377), .A2(n724), .B0(n782), .B1(n1153), .Y(
        n793) );
  MX2 U839 ( .A(n783), .B(n784), .S0(n1155), .Y(n794) );
  MX2 U840 ( .A(n785), .B(n786), .S0(n1156), .Y(n795) );
  MX2 U841 ( .A(n787), .B(n788), .S0(n1124), .Y(n796) );
  OAI32 U842 ( .A0(n1122), .A1(n789), .A2(n790), .B0(n1123), .B1(n791), .Y(
        n797) );
  MX2 U843 ( .A(n792), .B(n793), .S0(n1123), .Y(n798) );
  MX2 U844 ( .A(n794), .B(n795), .S0(n1124), .Y(n799) );
  MX2 U845 ( .A(n796), .B(n797), .S0(n1129), .Y(n800) );
  MX2 U846 ( .A(n798), .B(n799), .S0(n1126), .Y(n801) );
  MX2 U847 ( .A(n800), .B(n801), .S0(n1143), .Y(\r_p_r/N3459 ) );
  MX2 U848 ( .A(n697), .B(n687), .S0(n1143), .Y(n802) );
  MX2 U849 ( .A(n1386), .B(n713), .S0(n1096), .Y(n803) );
  MX2 U850 ( .A(n802), .B(n803), .S0(n1127), .Y(n804) );
  MX2 U851 ( .A(n1086), .B(n1105), .S0(n1144), .Y(n805) );
  MX2 U852 ( .A(n1385), .B(n1085), .S0(n1119), .Y(n806) );
  MX2 U853 ( .A(n1092), .B(n1105), .S0(n1095), .Y(n807) );
  MX2 U854 ( .A(n722), .B(n1382), .S0(n1095), .Y(n808) );
  MX2 U855 ( .A(n658), .B(n1369), .S0(n1128), .Y(n809) );
  AOI32 U856 ( .A0(n651), .A1(n1142), .A2(n716), .B0(n1143), .B1(n703), .Y(
        n810) );
  MX2 U857 ( .A(n1385), .B(n805), .S0(n711), .Y(n811) );
  AOI32 U858 ( .A0(n1383), .A1(n1142), .A2(n716), .B0(n1095), .B1(n1372), .Y(
        n812) );
  MX2 U859 ( .A(n1383), .B(n806), .S0(n1097), .Y(n813) );
  MX2 U860 ( .A(n707), .B(n719), .S0(n1143), .Y(n814) );
  MX2 U861 ( .A(n715), .B(n1120), .S0(\r_p_r/counter_r[4] ), .Y(n815) );
  MX2 U862 ( .A(n807), .B(n712), .S0(n1129), .Y(n816) );
  MX2 U863 ( .A(n677), .B(n808), .S0(n1126), .Y(n817) );
  NOR2B U864 ( .AN(n1142), .B(n809), .Y(n818) );
  MX2 U865 ( .A(n810), .B(n811), .S0(n1127), .Y(n819) );
  MX2 U866 ( .A(n723), .B(n1179), .S0(n1128), .Y(n820) );
  MX2 U867 ( .A(n1384), .B(n812), .S0(n1129), .Y(n821) );
  AOI21 U868 ( .A0(n1121), .A1(n1125), .B0(n1095), .Y(n822) );
  MX2 U869 ( .A(n657), .B(n1382), .S0(n1126), .Y(n823) );
  MX2 U870 ( .A(n1375), .B(n1158), .S0(n1127), .Y(n824) );
  MX2 U871 ( .A(n813), .B(n814), .S0(n1128), .Y(n825) );
  MX2 U872 ( .A(n721), .B(n815), .S0(n1129), .Y(n826) );
  MX2 U873 ( .A(n816), .B(n817), .S0(n1157), .Y(n827) );
  MX2 U874 ( .A(n818), .B(n819), .S0(n1155), .Y(n828) );
  MX2 U876 ( .A(n820), .B(n821), .S0(n1154), .Y(n830) );
  NOR2 U877 ( .A(n1096), .B(n1153), .Y(n831) );
  AOI32 U878 ( .A0(n822), .A1(n1153), .A2(n823), .B0(n1154), .B1(n824), .Y(
        n832) );
  MX2 U879 ( .A(n825), .B(n826), .S0(n1155), .Y(n833) );
  MX2 U880 ( .A(n827), .B(n828), .S0(n1123), .Y(n834) );
  MX2 U881 ( .A(n829), .B(n830), .S0(n1124), .Y(n835) );
  OAI32 U882 ( .A0(n1122), .A1(n831), .A2(n832), .B0(n1124), .B1(n833), .Y(
        n836) );
  MX2 U883 ( .A(n834), .B(n835), .S0(n1116), .Y(n837) );
  NOR2 U884 ( .A(n836), .B(n1117), .Y(n838) );
  MX2 U885 ( .A(n837), .B(n838), .S0(n1114), .Y(\r_p_r/N3460 ) );
  MX2 U886 ( .A(n1104), .B(n1086), .S0(n1120), .Y(n839) );
  NOR2B U887 ( .AN(n716), .B(n1158), .Y(n840) );
  MX2 U888 ( .A(n662), .B(n1383), .S0(n1121), .Y(n841) );
  MX2 U889 ( .A(n701), .B(n655), .S0(n1097), .Y(n842) );
  MX2 U890 ( .A(n1092), .B(n1158), .S0(n1096), .Y(n843) );
  MX2 U892 ( .A(n839), .B(n703), .S0(n1095), .Y(n845) );
  MX2 U893 ( .A(n1105), .B(n840), .S0(n1142), .Y(n846) );
  MX2 U894 ( .A(n1158), .B(n719), .S0(n1096), .Y(n847) );
  NOR2B U895 ( .AN(n718), .B(n1375), .Y(n848) );
  MX2 U896 ( .A(n1158), .B(n1119), .S0(n1144), .Y(n849) );
  MX2 U897 ( .A(n841), .B(n1099), .S0(n1097), .Y(n850) );
  NOR2 U898 ( .A(n1095), .B(n662), .Y(n851) );
  MX2 U899 ( .A(n1105), .B(n662), .S0(\r_p_r/counter_r[4] ), .Y(n852) );
  MX2 U900 ( .A(n673), .B(n712), .S0(n1126), .Y(n853) );
  MX2 U901 ( .A(n842), .B(n843), .S0(n1127), .Y(n854) );
  MX2 U902 ( .A(n659), .B(n710), .S0(n1128), .Y(n855) );
  AOI32 U903 ( .A0(n664), .A1(n1127), .A2(n844), .B0(n845), .B1(n1125), .Y(
        n856) );
  MX2 U905 ( .A(n715), .B(n1375), .S0(n1129), .Y(n858) );
  MX2 U906 ( .A(n671), .B(n846), .S0(n1126), .Y(n859) );
  MX2 U907 ( .A(n847), .B(n848), .S0(n1125), .Y(n860) );
  MX2 U908 ( .A(n721), .B(n849), .S0(n1127), .Y(n861) );
  MX2 U909 ( .A(n850), .B(n851), .S0(n1128), .Y(n862) );
  AOI32 U910 ( .A0(n717), .A1(n1125), .A2(n718), .B0(n1128), .B1(n852), .Y(
        n863) );
  MX2 U911 ( .A(n853), .B(n854), .S0(\r_p_r/counter_r[5] ), .Y(n864) );
  MX2 U912 ( .A(n855), .B(n856), .S0(n1154), .Y(n865) );
  MX2 U913 ( .A(n804), .B(n857), .S0(n1157), .Y(n866) );
  AOI32 U914 ( .A0(n1144), .A1(n1153), .A2(n858), .B0(n1154), .B1(n859), .Y(
        n867) );
  MX2 U915 ( .A(n860), .B(n861), .S0(n1154), .Y(n868) );
  MX2 U916 ( .A(n862), .B(n863), .S0(n1155), .Y(n869) );
  MX2 U917 ( .A(n864), .B(n865), .S0(n1123), .Y(n870) );
  MX2 U918 ( .A(n866), .B(n867), .S0(n1124), .Y(n871) );
  MX2 U919 ( .A(n868), .B(n869), .S0(n1123), .Y(n872) );
  MX2 U920 ( .A(n870), .B(n871), .S0(n1117), .Y(n873) );
  NOR2B U921 ( .AN(n872), .B(n1116), .Y(n874) );
  MX2 U922 ( .A(n873), .B(n874), .S0(n1113), .Y(\r_p_r/N3461 ) );
  NOR2 U923 ( .A(n1096), .B(n1104), .Y(n875) );
  MX2 U925 ( .A(n659), .B(n876), .S0(n1157), .Y(n877) );
  MX2 U926 ( .A(n693), .B(n665), .S0(n1144), .Y(n878) );
  NOR2B U927 ( .AN(n878), .B(n1153), .Y(n695) );
  NOR2 U928 ( .A(n1097), .B(n670), .Y(n879) );
  MX2 U930 ( .A(n1373), .B(n1386), .S0(n1144), .Y(n881) );
  MX2 U931 ( .A(n709), .B(n881), .S0(n1156), .Y(n882) );
  NOR2 U933 ( .A(n684), .B(n883), .Y(n884) );
  NOR2 U934 ( .A(n1143), .B(n1382), .Y(n885) );
  NOR2 U935 ( .A(n1367), .B(n1142), .Y(n886) );
  MX2 U936 ( .A(n651), .B(n1370), .S0(n1096), .Y(n887) );
  MX2 U937 ( .A(n1382), .B(n692), .S0(n1143), .Y(n888) );
  NOR2B U938 ( .AN(n710), .B(n1154), .Y(n889) );
  MX2 U939 ( .A(n675), .B(n660), .S0(n1143), .Y(n890) );
  MX2 U940 ( .A(n670), .B(n678), .S0(n1157), .Y(n891) );
  NOR2B U941 ( .AN(n880), .B(n884), .Y(n892) );
  MX2 U942 ( .A(n885), .B(n1098), .S0(n711), .Y(n893) );
  NOR2B U943 ( .AN(n681), .B(n705), .Y(n894) );
  AOI222 U944 ( .A0(n705), .A1(n1118), .B0(n705), .B1(n1382), .C0(n1118), .C1(
        n1143), .Y(n895) );
  NOR2B U945 ( .AN(n693), .B(n886), .Y(n896) );
  NOR2B U946 ( .AN(n690), .B(n1142), .Y(n897) );
  MX2 U947 ( .A(n1179), .B(n702), .S0(\r_p_r/counter_r[5] ), .Y(n898) );
  MX2 U948 ( .A(n887), .B(n888), .S0(n1156), .Y(n899) );
  OAI21 U950 ( .A0(n709), .A1(n1153), .B0(n698), .Y(n901) );
  MX2 U952 ( .A(n890), .B(n1371), .S0(n1155), .Y(n903) );
  MX2 U953 ( .A(n1104), .B(n891), .S0(n649), .Y(n904) );
  MX2 U954 ( .A(n892), .B(n893), .S0(n1156), .Y(n905) );
  MX2 U955 ( .A(n894), .B(n895), .S0(n1157), .Y(n906) );
  MX2 U956 ( .A(n896), .B(n897), .S0(n1155), .Y(n907) );
  MX2 U957 ( .A(n898), .B(n899), .S0(n1129), .Y(n908) );
  MX2 U958 ( .A(n877), .B(n900), .S0(n1126), .Y(n909) );
  MX2 U959 ( .A(n901), .B(n902), .S0(n1127), .Y(n910) );
  MX2 U960 ( .A(n903), .B(n904), .S0(n1128), .Y(n911) );
  MX2 U961 ( .A(n905), .B(n906), .S0(n1129), .Y(n912) );
  MX2 U962 ( .A(n907), .B(n882), .S0(n1126), .Y(n913) );
  MX2 U963 ( .A(n908), .B(n909), .S0(n1124), .Y(n914) );
  MX2 U964 ( .A(n910), .B(n911), .S0(n1123), .Y(n915) );
  MX2 U965 ( .A(n912), .B(n913), .S0(n1124), .Y(n916) );
  MX2 U966 ( .A(n914), .B(n915), .S0(n1116), .Y(n917) );
  NOR2B U967 ( .AN(n916), .B(n1117), .Y(n918) );
  MX2 U968 ( .A(n917), .B(n918), .S0(n1114), .Y(\r_p_r/N3462 ) );
  MX2 U969 ( .A(n665), .B(n666), .S0(n1143), .Y(n919) );
  MX2 U971 ( .A(n1382), .B(n1099), .S0(n1097), .Y(n920) );
  OAI221 U972 ( .A0(n1156), .A1(n700), .B0(n1153), .B1(n920), .C0(n1129), .Y(
        n921) );
  MX2 U973 ( .A(n1386), .B(n1099), .S0(n1144), .Y(n922) );
  MX2 U974 ( .A(n667), .B(n676), .S0(n1095), .Y(n923) );
  MX2 U975 ( .A(n922), .B(n923), .S0(n1154), .Y(n924) );
  NOR2B U976 ( .AN(n924), .B(n1126), .Y(n925) );
  MX2 U977 ( .A(n706), .B(n688), .S0(n1095), .Y(n926) );
  NOR2B U978 ( .AN(n926), .B(n1153), .Y(n927) );
  MX2 U979 ( .A(n657), .B(n662), .S0(n1119), .Y(n928) );
  MX2 U980 ( .A(n1382), .B(n1158), .S0(n1096), .Y(n929) );
  AOI221 U981 ( .A0(n701), .A1(n880), .B0(n1142), .B1(n880), .C0(n1156), .Y(
        n930) );
  MX2 U982 ( .A(n1158), .B(n1092), .S0(n1143), .Y(n931) );
  MX2 U983 ( .A(n1374), .B(n928), .S0(\r_p_r/counter_r[4] ), .Y(n932) );
  MX2 U984 ( .A(n1086), .B(n1385), .S0(n1120), .Y(n933) );
  MX2 U985 ( .A(n660), .B(n707), .S0(n1096), .Y(n934) );
  MX2 U986 ( .A(n929), .B(n661), .S0(n1155), .Y(n935) );
  OAI221 U988 ( .A0(n1157), .A1(n702), .B0(n1153), .B1(n679), .C0(n1127), .Y(
        n937) );
  NOR2 U989 ( .A(n927), .B(n930), .Y(n938) );
  MX2 U990 ( .A(n931), .B(n932), .S0(\r_p_r/counter_r[5] ), .Y(n939) );
  AOI32 U991 ( .A0(n1096), .A1(n1153), .A2(n933), .B0(n1157), .B1(n668), .Y(
        n940) );
  AOI32 U992 ( .A0(n1155), .A1(n1125), .A2(n934), .B0(n1128), .B1(n935), .Y(
        n941) );
  MX2 U993 ( .A(n877), .B(n694), .S0(n1127), .Y(n942) );
  AOI32 U994 ( .A0(n698), .A1(n921), .A2(n936), .B0(n1129), .B1(n921), .Y(n943) );
  MX2 U996 ( .A(n938), .B(n939), .S0(n1128), .Y(n945) );
  MX2 U997 ( .A(n940), .B(n882), .S0(n1129), .Y(n946) );
  MX2 U998 ( .A(n941), .B(n942), .S0(n1123), .Y(n947) );
  MX2 U999 ( .A(n943), .B(n944), .S0(n1124), .Y(n948) );
  MX2 U1000 ( .A(n945), .B(n946), .S0(n1123), .Y(n949) );
  MX2 U1001 ( .A(n947), .B(n948), .S0(n1117), .Y(n950) );
  NOR2B U1002 ( .AN(n949), .B(n1116), .Y(n951) );
  MX2 U1003 ( .A(n950), .B(n951), .S0(n1113), .Y(\r_p_r/N3463 ) );
  MX2 U1004 ( .A(n1375), .B(n682), .S0(n1097), .Y(n952) );
  NOR2B U1005 ( .AN(n952), .B(\r_p_r/counter_r[5] ), .Y(n953) );
  MX2 U1006 ( .A(n690), .B(n691), .S0(n1154), .Y(n954) );
  MX2 U1007 ( .A(n1386), .B(n1099), .S0(n1121), .Y(n955) );
  NOR2 U1008 ( .A(n1096), .B(n1375), .Y(n956) );
  NOR2 U1010 ( .A(n954), .B(n649), .Y(n958) );
  MX2 U1011 ( .A(n1105), .B(n955), .S0(n1095), .Y(n959) );
  MX2 U1012 ( .A(n678), .B(n1098), .S0(n1095), .Y(n960) );
  NOR2 U1013 ( .A(n1156), .B(n956), .Y(n961) );
  MX2 U1014 ( .A(n1385), .B(n1092), .S0(n1095), .Y(n962) );
  MX2 U1015 ( .A(n663), .B(n1372), .S0(n1096), .Y(n963) );
  MX2 U1016 ( .A(n957), .B(n1373), .S0(\r_p_r/counter_r[4] ), .Y(n964) );
  MX2 U1017 ( .A(n958), .B(n692), .S0(n1126), .Y(n965) );
  NOR2B U1018 ( .AN(n1126), .B(n1159), .Y(n966) );
  MX2 U1019 ( .A(n659), .B(n959), .S0(n1157), .Y(n967) );
  AOI221 U1020 ( .A0(n1143), .A1(n698), .B0(n699), .B1(n698), .C0(n1127), .Y(
        n968) );
  OAI221 U1021 ( .A0(n1156), .A1(n702), .B0(n1153), .B1(n960), .C0(n1128), .Y(
        n969) );
  NOR2 U1022 ( .A(n961), .B(n927), .Y(n970) );
  MX2 U1023 ( .A(n962), .B(n689), .S0(n1154), .Y(n971) );
  AOI221 U1024 ( .A0(n704), .A1(n1154), .B0(n705), .B1(n1157), .C0(n953), .Y(
        n972) );
  MX2 U1025 ( .A(n963), .B(n964), .S0(n1155), .Y(n973) );
  NOR2B U1026 ( .AN(n965), .B(n966), .Y(n974) );
  MX2 U1027 ( .A(n967), .B(n694), .S0(n1127), .Y(n975) );
  MX2 U1030 ( .A(n970), .B(n971), .S0(n1128), .Y(n978) );
  MX2 U1031 ( .A(n972), .B(n973), .S0(n1129), .Y(n979) );
  MX2 U1032 ( .A(n974), .B(n975), .S0(n1124), .Y(n980) );
  MX2 U1033 ( .A(n976), .B(n977), .S0(n1123), .Y(n981) );
  MX2 U1034 ( .A(n978), .B(n979), .S0(n1124), .Y(n982) );
  MX2 U1035 ( .A(n980), .B(n981), .S0(n1116), .Y(n983) );
  NOR2B U1036 ( .AN(n982), .B(n1117), .Y(n984) );
  MX2 U1037 ( .A(n983), .B(n984), .S0(n1114), .Y(\r_p_r/N3464 ) );
  MX2 U1038 ( .A(n1092), .B(n1158), .S0(n1157), .Y(n985) );
  MX2 U1039 ( .A(n1099), .B(n1158), .S0(n1119), .Y(n986) );
  MX2 U1040 ( .A(n1382), .B(n1386), .S0(n1120), .Y(n987) );
  NOR2B U1041 ( .AN(n985), .B(n649), .Y(n988) );
  MX2 U1042 ( .A(n669), .B(n670), .S0(n1144), .Y(n989) );
  MX2 U1043 ( .A(n674), .B(n675), .S0(n1144), .Y(n990) );
  MX2 U1044 ( .A(n986), .B(n1383), .S0(n1097), .Y(n991) );
  MX2 U1045 ( .A(n655), .B(n987), .S0(n1144), .Y(n992) );
  MX2 U1046 ( .A(n686), .B(n1367), .S0(n1143), .Y(n993) );
  MX2 U1047 ( .A(n1375), .B(n1092), .S0(n1143), .Y(n994) );
  MX2 U1048 ( .A(n683), .B(n655), .S0(n1096), .Y(n995) );
  MX2 U1049 ( .A(n685), .B(n1104), .S0(n1144), .Y(n996) );
  MX2 U1050 ( .A(n655), .B(n988), .S0(n1126), .Y(n997) );
  NOR2 U1051 ( .A(n1129), .B(n1159), .Y(n998) );
  MX2 U1052 ( .A(n659), .B(n661), .S0(n1156), .Y(n999) );
  AOI32 U1053 ( .A0(n664), .A1(n696), .A2(n668), .B0(n1153), .B1(n696), .Y(
        n1000) );
  MX2 U1054 ( .A(n989), .B(n671), .S0(n1157), .Y(n1001) );
  MX2 U1055 ( .A(n672), .B(n673), .S0(\r_p_r/counter_r[5] ), .Y(n1002) );
  MX2 U1056 ( .A(n990), .B(n991), .S0(n1156), .Y(n1003) );
  MX2 U1057 ( .A(n677), .B(n679), .S0(n1155), .Y(n1004) );
  MX2 U1058 ( .A(n992), .B(n993), .S0(n1156), .Y(n1005) );
  MX2 U1059 ( .A(n994), .B(n689), .S0(n1156), .Y(n1006) );
  AOI221 U1060 ( .A0(n670), .A1(n1155), .B0(n681), .B1(n1155), .C0(n953), .Y(
        n1007) );
  MX2 U1061 ( .A(n995), .B(n996), .S0(n1155), .Y(n1008) );
  NOR2B U1062 ( .AN(n997), .B(n998), .Y(n1009) );
  MX2 U1063 ( .A(n999), .B(n1000), .S0(n1127), .Y(n1010) );
  MX2 U1064 ( .A(n1001), .B(n1002), .S0(n1128), .Y(n1011) );
  MX2 U1065 ( .A(n1003), .B(n1004), .S0(n1129), .Y(n1012) );
  MX2 U1066 ( .A(n1005), .B(n1006), .S0(n1126), .Y(n1013) );
  MX2 U1067 ( .A(n1007), .B(n1008), .S0(n1127), .Y(n1014) );
  MX2 U1068 ( .A(n1009), .B(n1010), .S0(n1123), .Y(n1015) );
  MX2 U1069 ( .A(n1011), .B(n1012), .S0(n1124), .Y(n1016) );
  MX2 U1070 ( .A(n1013), .B(n1014), .S0(n1123), .Y(n1017) );
  MX2 U1071 ( .A(n1015), .B(n1016), .S0(n1117), .Y(n1018) );
  NOR2B U1072 ( .AN(n1017), .B(n1116), .Y(n1019) );
  MX2 U1073 ( .A(n1018), .B(n1019), .S0(n1113), .Y(\r_p_r/N3465 ) );
  MX2 U1074 ( .A(n714), .B(n1365), .S0(n1154), .Y(n1020) );
  MX2 U1076 ( .A(n1020), .B(n1160), .S0(n1128), .Y(n1022) );
  MX2 U1077 ( .A(n1368), .B(n1375), .S0(n1095), .Y(n1023) );
  MX2 U1078 ( .A(n1105), .B(n708), .S0(n1095), .Y(n1024) );
  MX2 U1079 ( .A(n1023), .B(n1024), .S0(n1155), .Y(n1025) );
  AND2 U1080 ( .A(n1095), .B(n666), .Y(n1026) );
  MX2 U1082 ( .A(n693), .B(n667), .S0(n1097), .Y(n1028) );
  MX2 U1083 ( .A(n1027), .B(n1028), .S0(\r_p_r/counter_r[5] ), .Y(n1029) );
  MX2 U1084 ( .A(n1025), .B(n1029), .S0(n1129), .Y(n1030) );
  MX2 U1085 ( .A(n1022), .B(n1030), .S0(n1124), .Y(n1031) );
  AOI2BB1 U1086 ( .A0N(n1142), .A1N(n683), .B0(n1372), .Y(n1032) );
  MX2 U1087 ( .A(n1098), .B(n1086), .S0(n1121), .Y(n1033) );
  MX2 U1088 ( .A(n1377), .B(n1033), .S0(n1143), .Y(n1034) );
  MX2 U1089 ( .A(n1032), .B(n1034), .S0(n1154), .Y(n1035) );
  NOR2B U1090 ( .AN(n693), .B(n683), .Y(n1036) );
  NOR2B U1091 ( .AN(n1367), .B(n1382), .Y(n1037) );
  MX2 U1092 ( .A(n1036), .B(n1037), .S0(\r_p_r/counter_r[4] ), .Y(n1038) );
  NOR2B U1093 ( .AN(n1038), .B(n1153), .Y(n1039) );
  MX2 U1094 ( .A(n1035), .B(n1039), .S0(n1126), .Y(n1040) );
  MX2 U1095 ( .A(n674), .B(n1383), .S0(n1095), .Y(n1041) );
  MX2 U1096 ( .A(n1380), .B(n708), .S0(n1096), .Y(n1042) );
  MX2 U1097 ( .A(n1041), .B(n1042), .S0(n1157), .Y(n1043) );
  MX2 U1099 ( .A(n680), .B(n707), .S0(n1144), .Y(n1045) );
  AOI221 U1100 ( .A0(n1044), .A1(n1157), .B0(n1144), .B1(n1154), .C0(n1045), 
        .Y(n1046) );
  MX2 U1101 ( .A(n1043), .B(n1046), .S0(n1127), .Y(n1047) );
  MX2 U1102 ( .A(n1040), .B(n1047), .S0(n1123), .Y(n1048) );
  MX2 U1103 ( .A(n1031), .B(n1048), .S0(n1116), .Y(n1049) );
  MX2 U1104 ( .A(n655), .B(n651), .S0(n1144), .Y(n1050) );
  NOR2B U1105 ( .AN(n686), .B(n1092), .Y(n1051) );
  MX2 U1106 ( .A(n1367), .B(n1051), .S0(n1142), .Y(n1052) );
  MX2 U1107 ( .A(n1050), .B(n1052), .S0(n1154), .Y(n1053) );
  AOI32 U1109 ( .A0(n1142), .A1(n1378), .A2(n657), .B0(n719), .B1(n1097), .Y(
        n1055) );
  MX2 U1110 ( .A(n1054), .B(n1055), .S0(n1156), .Y(n1056) );
  MX2 U1111 ( .A(n1053), .B(n1056), .S0(n1128), .Y(n1057) );
  MX2 U1112 ( .A(n685), .B(n1376), .S0(n1096), .Y(n1058) );
  NOR2B U1113 ( .AN(n707), .B(n1142), .Y(n1059) );
  MX2 U1114 ( .A(n1058), .B(n1059), .S0(n1157), .Y(n1060) );
  MX2 U1115 ( .A(n663), .B(n688), .S0(n1097), .Y(n1061) );
  MX2 U1116 ( .A(n1370), .B(n1104), .S0(n1095), .Y(n1062) );
  MX2 U1117 ( .A(n1061), .B(n1062), .S0(n1156), .Y(n1063) );
  MX2 U1118 ( .A(n1060), .B(n1063), .S0(n1129), .Y(n1064) );
  MX2 U1119 ( .A(n1057), .B(n1064), .S0(n1124), .Y(n1065) );
  NOR2B U1120 ( .AN(n1065), .B(n1117), .Y(n1066) );
  MX2 U1121 ( .A(n1049), .B(n1066), .S0(n1114), .Y(\r_p_r/N3466 ) );
  OR2 U1128 ( .A(n1137), .B(n1402), .Y(n1073) );
  OR2 U1129 ( .A(n1137), .B(n211), .Y(n1074) );
  OR2 U1130 ( .A(n1135), .B(n1398), .Y(n1075) );
  OR2 U1131 ( .A(n1119), .B(n651), .Y(n1076) );
  OR2 U1132 ( .A(n1137), .B(n1163), .Y(n1077) );
  INV U1133 ( .A(n228), .Y(n1078) );
  INV U1134 ( .A(n1078), .Y(n1079) );
  INV U1135 ( .A(n1075), .Y(n1080) );
  INV U1136 ( .A(n1073), .Y(n1081) );
  INV U1137 ( .A(n1074), .Y(n1082) );
  INV U1138 ( .A(n227), .Y(n1083) );
  INV U1139 ( .A(n1083), .Y(n1084) );
  INV U1140 ( .A(\r_p_r/counter_r[2] ), .Y(n1085) );
  INV U1141 ( .A(n1085), .Y(n1086) );
  INV U1142 ( .A(n232), .Y(n1087) );
  INV U1143 ( .A(n1087), .Y(n1088) );
  INV U1144 ( .A(n1077), .Y(n1089) );
  INV U1145 ( .A(n1149), .Y(n1090) );
  INV U1146 ( .A(n1149), .Y(n1091) );
  INV U1147 ( .A(n1076), .Y(n1092) );
  INV U1148 ( .A(n1145), .Y(n1093) );
  INV U1149 ( .A(n1145), .Y(n1094) );
  INV U1150 ( .A(n1142), .Y(n1095) );
  INV U1151 ( .A(n1142), .Y(n1096) );
  INV U1152 ( .A(n1142), .Y(n1097) );
  INV U1153 ( .A(n654), .Y(n1098) );
  INV U1154 ( .A(n1098), .Y(n1099) );
  INV U1155 ( .A(\l_p_r/counter_r[0] ), .Y(n1100) );
  INV U1156 ( .A(n1100), .Y(n1101) );
  INV U1157 ( .A(\l_p_r/counter_r[1] ), .Y(n1102) );
  INV U1158 ( .A(n1102), .Y(n1103) );
  INV U1159 ( .A(\r_p_r/counter_r[3] ), .Y(n1104) );
  INV U1160 ( .A(n1104), .Y(n1105) );
  INV U1161 ( .A(\l_p_r/counter_r[6] ), .Y(n1106) );
  INV U1162 ( .A(n1106), .Y(n1107) );
  INV U1163 ( .A(n1106), .Y(n1108) );
  INV U1164 ( .A(\l_p_r/counter_r[7] ), .Y(n1109) );
  INV U1165 ( .A(n1109), .Y(n1110) );
  INV U1166 ( .A(n1109), .Y(n1111) );
  INV U1167 ( .A(\r_p_r/counter_r[8] ), .Y(n1112) );
  INV U1168 ( .A(n1112), .Y(n1113) );
  INV U1169 ( .A(n1112), .Y(n1114) );
  INV U1170 ( .A(\r_p_r/counter_r[7] ), .Y(n1115) );
  INV U1171 ( .A(n1115), .Y(n1116) );
  INV U1172 ( .A(n1115), .Y(n1117) );
  INV U1173 ( .A(\r_p_r/counter_r[0] ), .Y(n1118) );
  INV U1174 ( .A(n1118), .Y(n1119) );
  INV U1175 ( .A(n1118), .Y(n1120) );
  INV U1176 ( .A(n1118), .Y(n1121) );
  INV U1177 ( .A(\r_p_r/counter_r[6] ), .Y(n1122) );
  INV U1178 ( .A(n1122), .Y(n1123) );
  INV U1179 ( .A(n1122), .Y(n1124) );
  INV U1180 ( .A(\r_p_r/counter_r[1] ), .Y(n1125) );
  INV U1181 ( .A(n1125), .Y(n1126) );
  INV U1182 ( .A(n1125), .Y(n1127) );
  INV U1183 ( .A(n1125), .Y(n1128) );
  INV U1184 ( .A(n1125), .Y(n1129) );
  INV U1185 ( .A(\l_p_r/counter_r[8] ), .Y(n1130) );
  INV U1186 ( .A(n1130), .Y(n1131) );
  INV U1187 ( .A(n1130), .Y(n1132) );
  INV U1188 ( .A(n1130), .Y(n1133) );
  INV U1189 ( .A(\l_p_r/counter_r[5] ), .Y(n1134) );
  INV U1190 ( .A(n1134), .Y(n1135) );
  INV U1191 ( .A(n1134), .Y(n1136) );
  INV U1192 ( .A(n1134), .Y(n1137) );
  INV U1193 ( .A(\l_p_r/counter_r[4] ), .Y(n1138) );
  INV U1194 ( .A(n1138), .Y(n1139) );
  INV U1195 ( .A(n1138), .Y(n1140) );
  INV U1196 ( .A(n1138), .Y(n1141) );
  INV U1197 ( .A(\r_p_r/counter_r[4] ), .Y(n1142) );
  INV U1198 ( .A(n1142), .Y(n1143) );
  INV U1199 ( .A(n1142), .Y(n1144) );
  INV U1200 ( .A(\l_p_r/counter_r[3] ), .Y(n1145) );
  INV U1201 ( .A(n1145), .Y(n1146) );
  INV U1202 ( .A(n1145), .Y(n1147) );
  INV U1203 ( .A(n1145), .Y(n1148) );
  INV U1204 ( .A(\l_p_r/counter_r[2] ), .Y(n1149) );
  INV U1205 ( .A(n1149), .Y(n1150) );
  INV U1206 ( .A(n1149), .Y(n1151) );
  INV U1207 ( .A(n1149), .Y(n1152) );
  INV U1208 ( .A(\r_p_r/counter_r[5] ), .Y(n1153) );
  INV U1209 ( .A(n1153), .Y(n1154) );
  INV U1210 ( .A(n1153), .Y(n1155) );
  INV U1211 ( .A(n1153), .Y(n1156) );
  INV U1212 ( .A(n1153), .Y(n1157) );
  AND2 U1213 ( .A(n1086), .B(n1105), .Y(n1158) );
  AND2 U1214 ( .A(n1144), .B(n1155), .Y(n1159) );
  AND2 U1215 ( .A(n692), .B(n1159), .Y(n1160) );
  AND2 U1216 ( .A(n235), .B(n215), .Y(n1161) );
  AND2 U1217 ( .A(n230), .B(n235), .Y(n1162) );
  LOGIC_0 U1218 ( .LOGIC_0_PIN(\g_l_d1/*Logic0* ) );
  INV U1219 ( .A(\l_p_r/N2849 ), .Y(n1339) );
  OAI22 U1220 ( .A0(n1133), .A1(graphic_lcd_en), .B0(n1301), .B1(
        graphic_lcd_en), .Y(n1300) );
  INV U1221 ( .A(n1220), .Y(n1212) );
  INV U1222 ( .A(\r_p_r/N3458 ), .Y(n1340) );
  OAI21 U1223 ( .A0(graphic_lcd_en), .A1(n1333), .B0(n1332), .Y(n1307) );
  NAND2B U1224 ( .AN(n1103), .B(n1101), .Y(n208) );
  NAND2B U1225 ( .AN(n214), .B(n1137), .Y(n215) );
  NAND2B U1226 ( .AN(n211), .B(n1135), .Y(n230) );
  NAND2B U1227 ( .AN(n1136), .B(n208), .Y(n235) );
  NAND2B U1228 ( .AN(n1392), .B(n1137), .Y(n236) );
  NAND2B U1229 ( .AN(n1135), .B(n1163), .Y(n237) );
  INV U1230 ( .A(n223), .Y(n1163) );
  NAND2B U1231 ( .AN(n1402), .B(n1136), .Y(n240) );
  NAND2B U1232 ( .AN(n220), .B(n1077), .Y(n251) );
  NAND2B U1233 ( .AN(n1134), .B(n1392), .Y(n258) );
  NAND2B U1234 ( .AN(n212), .B(n1073), .Y(n262) );
  NAND2B U1235 ( .AN(n1088), .B(n258), .Y(n266) );
  NAND2B U1236 ( .AN(n1132), .B(n268), .Y(n269) );
  NAND2B U1237 ( .AN(n1133), .B(n263), .Y(n274) );
  NAND2B U1238 ( .AN(n1409), .B(n213), .Y(n277) );
  NAND2B U1239 ( .AN(n223), .B(n230), .Y(n279) );
  NAND2B U1240 ( .AN(n1134), .B(n1101), .Y(n280) );
  NAND2B U1241 ( .AN(n1131), .B(n1084), .Y(n288) );
  NAND2B U1242 ( .AN(n301), .B(n302), .Y(\l_p_r/N2849 ) );
  NAND2B U1243 ( .AN(n1148), .B(n1149), .Y(n332) );
  NAND2B U1244 ( .AN(n1084), .B(n1073), .Y(n344) );
  NAND2B U1245 ( .AN(n264), .B(n1164), .Y(n354) );
  INV U1246 ( .A(n352), .Y(n1164) );
  NAND2B U1247 ( .AN(n242), .B(n1111), .Y(n458) );
  NAND2B U1248 ( .AN(n1108), .B(n1132), .Y(n477) );
  NAND2B U1249 ( .AN(n1411), .B(n1150), .Y(n512) );
  NAND2B U1250 ( .AN(n1133), .B(n1165), .Y(n556) );
  INV U1251 ( .A(n546), .Y(n1165) );
  NAND2B U1252 ( .AN(n1147), .B(n237), .Y(n576) );
  NAND2B U1253 ( .AN(n1105), .B(n1085), .Y(n651) );
  NAND2B U1254 ( .AN(n656), .B(n657), .Y(n658) );
  NAND2B U1255 ( .AN(n1105), .B(n1086), .Y(n662) );
  NAND2B U1256 ( .AN(n1144), .B(n1166), .Y(n664) );
  INV U1257 ( .A(n663), .Y(n1166) );
  NAND2B U1258 ( .AN(n1120), .B(n651), .Y(n666) );
  NAND2B U1259 ( .AN(n1142), .B(n667), .Y(n668) );
  NAND2B U1260 ( .AN(n1121), .B(n1158), .Y(n676) );
  NAND2B U1261 ( .AN(n680), .B(n1143), .Y(n681) );
  NAND2B U1262 ( .AN(n1382), .B(n1167), .Y(n685) );
  INV U1263 ( .A(n684), .Y(n1167) );
  NAND2B U1264 ( .AN(n1385), .B(n1119), .Y(n686) );
  NAND2B U1265 ( .AN(n1099), .B(n1378), .Y(n688) );
  NAND2B U1266 ( .AN(n1118), .B(n1105), .Y(n691) );
  NAND2B U1267 ( .AN(n1120), .B(n1086), .Y(n693) );
  NAND2B U1268 ( .AN(n695), .B(n696), .Y(n694) );
  NAND2B U1269 ( .AN(n1153), .B(n685), .Y(n699) );
  NAND2B U1270 ( .AN(n657), .B(n1121), .Y(n716) );
  NAND2B U1271 ( .AN(n1119), .B(n1099), .Y(n717) );
  NAND2B U1272 ( .AN(n706), .B(n1096), .Y(n718) );
  NAND2B U1273 ( .AN(n1142), .B(n1366), .Y(n723) );
  NAND2B U1274 ( .AN(n1114), .B(n1116), .Y(n724) );
  NAND2B U1275 ( .AN(n1113), .B(n1386), .Y(n725) );
  NAND2B U1276 ( .AN(n1115), .B(n1154), .Y(n729) );
  NAND2B U1277 ( .AN(n747), .B(n748), .Y(\r_p_r/N3458 ) );
  NAND2B U1278 ( .AN(n1114), .B(n1168), .Y(n760) );
  INV U1279 ( .A(n722), .Y(n1168) );
  NAND2B U1280 ( .AN(n1113), .B(n1169), .Y(n765) );
  INV U1281 ( .A(n680), .Y(n1169) );
  NAND2B U1282 ( .AN(n1154), .B(n1170), .Y(n829) );
  INV U1283 ( .A(n804), .Y(n1170) );
  NAND2B U1284 ( .AN(n1142), .B(n665), .Y(n844) );
  NAND2B U1285 ( .AN(n1125), .B(n714), .Y(n857) );
  NAND2B U1286 ( .AN(n875), .B(n1171), .Y(n876) );
  INV U1287 ( .A(n704), .Y(n1171) );
  NAND2B U1288 ( .AN(n1386), .B(n879), .Y(n880) );
  NAND2B U1289 ( .AN(n1375), .B(n1097), .Y(n883) );
  NAND2B U1290 ( .AN(n695), .B(n1172), .Y(n900) );
  INV U1291 ( .A(n889), .Y(n1172) );
  NAND2B U1292 ( .AN(n1155), .B(n1173), .Y(n902) );
  INV U1293 ( .A(n700), .Y(n1173) );
  NAND2B U1294 ( .AN(n1154), .B(n919), .Y(n696) );
  OAI21 U1295 ( .A0(n708), .A1(n1142), .B0(n1174), .Y(n936) );
  INV U1296 ( .A(n699), .Y(n1174) );
  NAND2B U1297 ( .AN(n925), .B(n937), .Y(n944) );
  NAND2B U1298 ( .AN(n1120), .B(n1383), .Y(n957) );
  NAND2B U1299 ( .AN(n968), .B(n921), .Y(n976) );
  NAND2B U1300 ( .AN(n925), .B(n969), .Y(n977) );
  NAND2B U1301 ( .AN(n1026), .B(n880), .Y(n1027) );
  NAND2B U1302 ( .AN(n1105), .B(n1121), .Y(n1044) );
  NAND2B U1303 ( .AN(n1143), .B(n1175), .Y(n1054) );
  INV U1304 ( .A(n692), .Y(n1175) );
  NAND2 U1305 ( .A(n1101), .B(n1103), .Y(n1176) );
  INV U1306 ( .A(n1176), .Y(n211) );
  NAND2 U1307 ( .A(n211), .B(n1137), .Y(n1177) );
  INV U1308 ( .A(n1177), .Y(n212) );
  NAND2 U1309 ( .A(n1103), .B(n1135), .Y(n1178) );
  INV U1310 ( .A(n1178), .Y(n213) );
  NAND2 U1311 ( .A(n1158), .B(n1095), .Y(n1179) );
  INV U1312 ( .A(n1179), .Y(n672) );
  NAND2 U1313 ( .A(n1158), .B(n1119), .Y(n1180) );
  INV U1314 ( .A(n1180), .Y(n715) );
  NOR2 U1315 ( .A(n1181), .B(n1182), .Y(n1341) );
  XNOR2 U1316 ( .A(refresh), .B(n1183), .Y(n1181) );
  NOR2B U1317 ( .AN(\clk_div1/counter [13]), .B(n1184), .Y(n1183) );
  NOR2 U1318 ( .A(n1182), .B(n1185), .Y(n1342) );
  XOR2 U1319 ( .A(\clk_div1/counter [13]), .B(n1184), .Y(n1185) );
  NAND2 U1320 ( .A(n1186), .B(\clk_div1/counter [12]), .Y(n1184) );
  NOR2 U1321 ( .A(n1182), .B(n1187), .Y(n1343) );
  XNOR2 U1322 ( .A(n1186), .B(\clk_div1/counter [12]), .Y(n1187) );
  NOR2B U1323 ( .AN(\clk_div1/counter [11]), .B(n1188), .Y(n1186) );
  NOR2 U1324 ( .A(n1182), .B(n1189), .Y(n1344) );
  XOR2 U1325 ( .A(\clk_div1/counter [11]), .B(n1188), .Y(n1189) );
  NAND2 U1326 ( .A(n1190), .B(\clk_div1/counter [10]), .Y(n1188) );
  NOR2 U1327 ( .A(n1182), .B(n1191), .Y(n1345) );
  XNOR2 U1328 ( .A(n1190), .B(\clk_div1/counter [10]), .Y(n1191) );
  NOR2B U1329 ( .AN(\clk_div1/counter [9]), .B(n1192), .Y(n1190) );
  NOR2 U1330 ( .A(n1182), .B(n1193), .Y(n1346) );
  XOR2 U1331 ( .A(\clk_div1/counter [9]), .B(n1192), .Y(n1193) );
  NAND2 U1332 ( .A(n1194), .B(\clk_div1/counter [8]), .Y(n1192) );
  NOR2 U1333 ( .A(n1182), .B(n1195), .Y(n1347) );
  XNOR2 U1334 ( .A(n1194), .B(\clk_div1/counter [8]), .Y(n1195) );
  NOR2B U1335 ( .AN(\clk_div1/counter [7]), .B(n1196), .Y(n1194) );
  NOR2 U1336 ( .A(n1182), .B(n1197), .Y(n1348) );
  XOR2 U1337 ( .A(\clk_div1/counter [7]), .B(n1196), .Y(n1197) );
  NAND2 U1338 ( .A(n1198), .B(\clk_div1/counter [6]), .Y(n1196) );
  NOR2 U1339 ( .A(n1182), .B(n1199), .Y(n1349) );
  XNOR2 U1340 ( .A(n1198), .B(\clk_div1/counter [6]), .Y(n1199) );
  NOR2B U1341 ( .AN(\clk_div1/counter [5]), .B(n1200), .Y(n1198) );
  NOR2 U1342 ( .A(n1182), .B(n1201), .Y(n1350) );
  XOR2 U1343 ( .A(\clk_div1/counter [5]), .B(n1200), .Y(n1201) );
  NAND2 U1344 ( .A(n1202), .B(\clk_div1/counter [4]), .Y(n1200) );
  NOR2 U1345 ( .A(n1182), .B(n1203), .Y(n1351) );
  XNOR2 U1346 ( .A(n1202), .B(\clk_div1/counter [4]), .Y(n1203) );
  NOR2B U1347 ( .AN(\clk_div1/counter [3]), .B(n1204), .Y(n1202) );
  NOR2 U1348 ( .A(n1182), .B(n1205), .Y(n1352) );
  XOR2 U1349 ( .A(\clk_div1/counter [3]), .B(n1204), .Y(n1205) );
  NAND3 U1350 ( .A(\clk_div1/counter [2]), .B(\clk_div1/counter [0]), .C(
        \clk_div1/counter [1]), .Y(n1204) );
  OAI2BB2 U1351 ( .B0(n1206), .B1(n1207), .A0N(auto_i), .A1N(n1208), .Y(n1353)
         );
  MX2 U1352 ( .A(\clk_div1/counter [2]), .B(n1209), .S0(\clk_div1/counter [1]), 
        .Y(n1208) );
  NOR2B U1353 ( .AN(\clk_div1/counter [0]), .B(\clk_div1/counter [2]), .Y(
        n1209) );
  INV U1354 ( .A(n1355), .Y(n1207) );
  INV U1355 ( .A(\clk_div1/counter [2]), .Y(n1206) );
  MX2 U1356 ( .A(n1210), .B(n1355), .S0(\clk_div1/counter [1]), .Y(n1354) );
  NOR2B U1357 ( .AN(\clk_div1/counter [0]), .B(n1182), .Y(n1210) );
  INV U1358 ( .A(auto_i), .Y(n1182) );
  NOR2B U1359 ( .AN(auto_i), .B(\clk_div1/counter [0]), .Y(n1355) );
  INV U1360 ( .A(n1211), .Y(graphic_lcd_d[7]) );
  AOI22 U1361 ( .A0(n1212), .A1(\l_p_r/N2857 ), .B0(n1220), .B1(\r_p_r/N3466 ), 
        .Y(n1211) );
  INV U1362 ( .A(n1213), .Y(graphic_lcd_d[6]) );
  AOI22 U1363 ( .A0(n1212), .A1(\l_p_r/N2856 ), .B0(n1220), .B1(\r_p_r/N3465 ), 
        .Y(n1213) );
  INV U1364 ( .A(n1214), .Y(graphic_lcd_d[5]) );
  AOI22 U1365 ( .A0(n1212), .A1(\l_p_r/N2855 ), .B0(n1220), .B1(\r_p_r/N3464 ), 
        .Y(n1214) );
  INV U1366 ( .A(n1215), .Y(graphic_lcd_d[4]) );
  AOI22 U1367 ( .A0(n1212), .A1(\l_p_r/N2854 ), .B0(n1220), .B1(\r_p_r/N3463 ), 
        .Y(n1215) );
  INV U1368 ( .A(n1216), .Y(graphic_lcd_d[3]) );
  AOI22 U1369 ( .A0(n1212), .A1(\l_p_r/N2853 ), .B0(n1220), .B1(\r_p_r/N3462 ), 
        .Y(n1216) );
  INV U1370 ( .A(n1217), .Y(graphic_lcd_d[2]) );
  AOI22 U1371 ( .A0(n1212), .A1(\l_p_r/N2852 ), .B0(n1220), .B1(\r_p_r/N3461 ), 
        .Y(n1217) );
  INV U1372 ( .A(n1218), .Y(graphic_lcd_d[1]) );
  AOI22 U1373 ( .A0(n1212), .A1(\l_p_r/N2851 ), .B0(n1220), .B1(\r_p_r/N3460 ), 
        .Y(n1218) );
  INV U1374 ( .A(n1219), .Y(graphic_lcd_d[0]) );
  AOI22 U1375 ( .A0(n1212), .A1(\l_p_r/N2850 ), .B0(n1220), .B1(\r_p_r/N3459 ), 
        .Y(n1219) );
  INV U1376 ( .A(n723), .Y(n1365) );
  INV U1377 ( .A(n691), .Y(n1366) );
  INV U1378 ( .A(n656), .Y(n1367) );
  INV U1379 ( .A(n658), .Y(n1368) );
  INV U1380 ( .A(n665), .Y(n1369) );
  INV U1381 ( .A(n667), .Y(n1370) );
  INV U1382 ( .A(n671), .Y(n1371) );
  INV U1383 ( .A(n669), .Y(n1372) );
  INV U1384 ( .A(n674), .Y(n1373) );
  INV U1385 ( .A(n675), .Y(n1374) );
  INV U1386 ( .A(n676), .Y(n1375) );
  INV U1387 ( .A(n682), .Y(n1376) );
  INV U1388 ( .A(n686), .Y(n1377) );
  INV U1389 ( .A(n687), .Y(n1378) );
  INV U1390 ( .A(n701), .Y(n1379) );
  INV U1391 ( .A(n717), .Y(n1380) );
  INV U1392 ( .A(n720), .Y(n1381) );
  INV U1393 ( .A(n651), .Y(n1382) );
  INV U1394 ( .A(n1158), .Y(n1383) );
  INV U1395 ( .A(n705), .Y(n1384) );
  INV U1396 ( .A(n657), .Y(n1385) );
  INV U1397 ( .A(n662), .Y(n1386) );
  INV U1398 ( .A(n233), .Y(n1387) );
  INV U1399 ( .A(n235), .Y(n1388) );
  INV U1400 ( .A(n241), .Y(n1389) );
  INV U1401 ( .A(n266), .Y(n1390) );
  INV U1402 ( .A(n258), .Y(n1391) );
  INV U1403 ( .A(n208), .Y(n1392) );
  INV U1404 ( .A(n239), .Y(n1393) );
  INV U1405 ( .A(n279), .Y(n1394) );
  INV U1406 ( .A(n265), .Y(n1395) );
  INV U1407 ( .A(n282), .Y(n1396) );
  INV U1408 ( .A(n253), .Y(n1397) );
  INV U1409 ( .A(n214), .Y(n1398) );
  INV U1410 ( .A(n215), .Y(n1399) );
  INV U1411 ( .A(n278), .Y(n1400) );
  INV U1412 ( .A(n240), .Y(n1401) );
  INV U1413 ( .A(n216), .Y(n1402) );
  INV U1414 ( .A(n225), .Y(n1403) );
  INV U1415 ( .A(n222), .Y(n1404) );
  INV U1416 ( .A(n237), .Y(n1405) );
  INV U1417 ( .A(n231), .Y(n1406) );
  INV U1418 ( .A(n277), .Y(n1407) );
  INV U1419 ( .A(n243), .Y(n1408) );
  INV U1420 ( .A(n273), .Y(n1409) );
  INV U1421 ( .A(n286), .Y(n1410) );
  XOR2 U1422 ( .A(mode), .B(n1221), .Y(n86) );
  NOR3B U1423 ( .AN(\g_l_d1/state[2] ), .B(\g_l_d1/state[1] ), .C(n1222), .Y(
        n1221) );
  INV U1424 ( .A(\g_l_d1/state[0] ), .Y(n1222) );
  OAI2BB1 U1425 ( .A0N(\g_l_d1/state[1] ), .A1N(n1223), .B0(n1224), .Y(n205)
         );
  AOI31 U1426 ( .A0(n1225), .A1(\re_detect1/sample_r[0] ), .A2(n1226), .B0(
        \g_l_d1/state[2] ), .Y(n1224) );
  INV U1427 ( .A(\re_detect1/sample_r[1] ), .Y(n1226) );
  MX2 U1428 ( .A(n1227), .B(n1228), .S0(graphic_lcd_en), .Y(n204) );
  NOR2B U1429 ( .AN(\g_l_d1/state[2] ), .B(n1225), .Y(n1228) );
  NOR2B U1430 ( .AN(n1229), .B(n1230), .Y(n203) );
  XNOR2 U1431 ( .A(\g_l_d1/counter[9] ), .B(n1231), .Y(n1230) );
  NOR2B U1432 ( .AN(\g_l_d1/counter[8] ), .B(n1232), .Y(n1231) );
  MX2 U1433 ( .A(n1233), .B(n1234), .S0(\g_l_d1/state[1] ), .Y(n202) );
  OAI21 U1434 ( .A0(\g_l_d1/state[0] ), .A1(n1223), .B0(n1235), .Y(n1234) );
  OAI211 U1435 ( .A0(\g_l_d1/counter[6] ), .A1(n1236), .B0(n1237), .C0(n1238), 
        .Y(n1223) );
  OAI2BB1 U1436 ( .A0N(n1239), .A1N(\g_l_d1/counter[2] ), .B0(
        \g_l_d1/counter[6] ), .Y(n1238) );
  NOR4BB U1437 ( .AN(n1240), .BN(n1241), .C(n1242), .D(n1243), .Y(n1237) );
  MX2 U1438 ( .A(rst_n), .B(n1244), .S0(\g_l_d1/counter[5] ), .Y(n1243) );
  XOR2 U1439 ( .A(rst_n), .B(\g_l_d1/counter[8] ), .Y(n1242) );
  NOR4 U1440 ( .A(\g_l_d1/counter[9] ), .B(\g_l_d1/counter[7] ), .C(
        \g_l_d1/counter[1] ), .D(n1245), .Y(n1241) );
  XOR2 U1441 ( .A(rst_n), .B(\g_l_d1/counter[0] ), .Y(n1245) );
  MX2 U1442 ( .A(n1244), .B(rst_n), .S0(\g_l_d1/counter[4] ), .Y(n1240) );
  NOR2 U1443 ( .A(n1239), .B(\g_l_d1/counter[2] ), .Y(n1236) );
  NOR2B U1444 ( .AN(rst_n), .B(n1246), .Y(n1239) );
  XOR2 U1445 ( .A(mode), .B(\g_l_d1/state[0] ), .Y(n1246) );
  NOR4BB U1446 ( .AN(\g_l_d1/state[0] ), .BN(\re_detect1/sample_r[0] ), .C(
        \g_l_d1/state[2] ), .D(\re_detect1/sample_r[1] ), .Y(n1233) );
  OAI2BB1 U1447 ( .A0N(\g_l_d1/state[1] ), .A1N(\g_l_d1/state[0] ), .B0(n1229), 
        .Y(n201) );
  NOR2B U1448 ( .AN(n1229), .B(n1247), .Y(n200) );
  XOR2 U1449 ( .A(\g_l_d1/counter[8] ), .B(n1232), .Y(n1247) );
  NAND2 U1450 ( .A(\g_l_d1/counter[7] ), .B(n1248), .Y(n1232) );
  NOR2B U1451 ( .AN(n1229), .B(n1249), .Y(n199) );
  XNOR2 U1452 ( .A(\g_l_d1/counter[7] ), .B(n1248), .Y(n1249) );
  NOR4BB U1453 ( .AN(n1250), .BN(\g_l_d1/counter[5] ), .C(n1251), .D(n1252), 
        .Y(n1248) );
  INV U1454 ( .A(\g_l_d1/counter[6] ), .Y(n1251) );
  NOR2B U1455 ( .AN(n1229), .B(n1253), .Y(n198) );
  XNOR2 U1456 ( .A(\g_l_d1/counter[6] ), .B(n1254), .Y(n1253) );
  NOR2B U1457 ( .AN(\g_l_d1/counter[5] ), .B(n1255), .Y(n1254) );
  NOR2B U1458 ( .AN(n1229), .B(n1256), .Y(n197) );
  XOR2 U1459 ( .A(\g_l_d1/counter[5] ), .B(n1255), .Y(n1256) );
  NAND2 U1460 ( .A(n1250), .B(graphic_lcd_en), .Y(n1255) );
  NOR3B U1461 ( .AN(\g_l_d1/counter[4] ), .B(n1244), .C(n1257), .Y(n1250) );
  NOR2B U1462 ( .AN(n1229), .B(n1258), .Y(n196) );
  XNOR2 U1463 ( .A(\g_l_d1/counter[4] ), .B(n1259), .Y(n1258) );
  NOR2B U1464 ( .AN(n1260), .B(n1244), .Y(n1259) );
  INV U1465 ( .A(\g_l_d1/counter[3] ), .Y(n1244) );
  NOR2B U1466 ( .AN(n1229), .B(n1261), .Y(n195) );
  XNOR2 U1467 ( .A(\g_l_d1/counter[3] ), .B(n1260), .Y(n1261) );
  NOR2 U1468 ( .A(n1257), .B(n1252), .Y(n1260) );
  INV U1469 ( .A(graphic_lcd_en), .Y(n1252) );
  NAND3 U1470 ( .A(\g_l_d1/counter[2] ), .B(\g_l_d1/counter[1] ), .C(
        \g_l_d1/counter[0] ), .Y(n1257) );
  NOR2B U1471 ( .AN(n1229), .B(n1262), .Y(n194) );
  XNOR2 U1472 ( .A(\g_l_d1/counter[2] ), .B(n1263), .Y(n1262) );
  NOR2B U1473 ( .AN(\g_l_d1/counter[1] ), .B(n1264), .Y(n1263) );
  NOR2B U1474 ( .AN(n1229), .B(n1265), .Y(n193) );
  XOR2 U1475 ( .A(\g_l_d1/counter[1] ), .B(n1264), .Y(n1265) );
  NAND2 U1476 ( .A(\g_l_d1/counter[0] ), .B(graphic_lcd_en), .Y(n1264) );
  NOR2B U1477 ( .AN(n1229), .B(n1266), .Y(n192) );
  XNOR2 U1478 ( .A(\g_l_d1/counter[0] ), .B(graphic_lcd_en), .Y(n1266) );
  NAND2B U1479 ( .AN(\g_l_d1/state[1] ), .B(n1267), .Y(n1229) );
  NAND2B U1480 ( .AN(n206), .B(n1268), .Y(n191) );
  MX2 U1481 ( .A(graphic_lcd_cs2), .B(\g_l_d1/state[0] ), .S0(n1227), .Y(n1268) );
  NOR2B U1482 ( .AN(\g_l_d1/state[1] ), .B(\g_l_d1/state[2] ), .Y(n1227) );
  NOR2B U1483 ( .AN(n1225), .B(n1235), .Y(n206) );
  NOR2 U1484 ( .A(\g_l_d1/state[1] ), .B(\g_l_d1/state[0] ), .Y(n1225) );
  MX2 U1485 ( .A(n1269), .B(n1270), .S0(\g_l_d1/state[1] ), .Y(n190) );
  NOR2B U1486 ( .AN(\g_l_d1/state[2] ), .B(n1271), .Y(n1270) );
  INV U1487 ( .A(n1267), .Y(n1269) );
  XNOR2 U1488 ( .A(\g_l_d1/state[0] ), .B(n1235), .Y(n1267) );
  INV U1489 ( .A(\g_l_d1/state[2] ), .Y(n1235) );
  MX2 U1490 ( .A(n1273), .B(n1274), .S0(n1101), .Y(n188) );
  MX2 U1491 ( .A(n1275), .B(n1276), .S0(n1103), .Y(n187) );
  NOR2B U1492 ( .AN(n1273), .B(n1100), .Y(n1275) );
  MX2 U1493 ( .A(n1277), .B(n1278), .S0(n1090), .Y(n186) );
  OAI21 U1494 ( .A0(n1103), .A1(n1279), .B0(n1280), .Y(n1278) );
  INV U1495 ( .A(n1276), .Y(n1280) );
  OAI21 U1496 ( .A0(n1101), .A1(n1279), .B0(n1281), .Y(n1276) );
  NOR3B U1497 ( .AN(n1273), .B(n1100), .C(n1102), .Y(n1277) );
  MX2 U1498 ( .A(n1282), .B(n1283), .S0(\l_p_r/counter_r[3] ), .Y(n185) );
  NOR2B U1499 ( .AN(n1273), .B(n1284), .Y(n1282) );
  MX2 U1500 ( .A(n1285), .B(n1286), .S0(n1139), .Y(n184) );
  OAI21 U1501 ( .A0(n1094), .A1(n1279), .B0(n1287), .Y(n1286) );
  INV U1502 ( .A(n1283), .Y(n1287) );
  OAI2BB1 U1503 ( .A0N(n1288), .A1N(n1284), .B0(n1281), .Y(n1283) );
  INV U1504 ( .A(n1279), .Y(n1288) );
  NOR3B U1505 ( .AN(n1273), .B(n1411), .C(n1284), .Y(n1285) );
  MX2 U1506 ( .A(n1289), .B(n1290), .S0(n1135), .Y(n183) );
  NOR2B U1507 ( .AN(n1291), .B(n1292), .Y(n1289) );
  MX2 U1508 ( .A(n1293), .B(n1294), .S0(n1107), .Y(n182) );
  OAI21 U1509 ( .A0(n1136), .A1(n1279), .B0(n1295), .Y(n1294) );
  INV U1510 ( .A(n1290), .Y(n1295) );
  OAI21 U1511 ( .A0(n1291), .A1(n1279), .B0(n1281), .Y(n1290) );
  INV U1512 ( .A(n1274), .Y(n1281) );
  NOR3B U1513 ( .AN(n1291), .B(n1134), .C(n1292), .Y(n1293) );
  MX2 U1514 ( .A(n1296), .B(n1297), .S0(n1110), .Y(n181) );
  INV U1515 ( .A(n1272), .Y(n1297) );
  NOR2B U1516 ( .AN(n1298), .B(n1292), .Y(n1296) );
  INV U1517 ( .A(n1273), .Y(n1292) );
  OAI2BB2 U1518 ( .B0(n1272), .B1(n1130), .A0N(n1273), .A1N(n1299), .Y(n180)
         );
  NOR2B U1519 ( .AN(n1298), .B(n1109), .Y(n1299) );
  NOR2 U1520 ( .A(n1274), .B(n1279), .Y(n1273) );
  AOI2BB1 U1521 ( .A0N(n1298), .A1N(n1279), .B0(n1274), .Y(n1272) );
  NOR2 U1522 ( .A(n1300), .B(n1279), .Y(n1274) );
  OAI31 U1523 ( .A0(n1411), .A1(n1134), .A2(n1302), .B0(n1303), .Y(n1301) );
  NOR2 U1524 ( .A(n1107), .B(n1111), .Y(n1303) );
  OAI31 U1525 ( .A0(n1101), .A1(n1103), .A2(n1152), .B0(n1141), .Y(n1302) );
  MX2 U1526 ( .A(sync_right), .B(graphic_lcd_rst), .S0(mode), .Y(n1279) );
  NOR3B U1527 ( .AN(n1291), .B(n1134), .C(n1106), .Y(n1298) );
  NOR3B U1528 ( .AN(n1139), .B(n1411), .C(n1284), .Y(n1291) );
  NAND3 U1529 ( .A(n1101), .B(n1103), .C(n1091), .Y(n1284) );
  INV U1530 ( .A(\l_p_r/counter_r[3] ), .Y(n1411) );
  MX2 U1531 ( .A(n1305), .B(n1306), .S0(n1119), .Y(n178) );
  INV U1532 ( .A(n1307), .Y(n1306) );
  MX2 U1533 ( .A(n1308), .B(n1309), .S0(n1126), .Y(n177) );
  NOR2B U1534 ( .AN(n1305), .B(n1118), .Y(n1308) );
  MX2 U1535 ( .A(n1310), .B(n1311), .S0(n1086), .Y(n176) );
  OAI21 U1536 ( .A0(n1127), .A1(n1312), .B0(n1313), .Y(n1311) );
  INV U1537 ( .A(n1309), .Y(n1313) );
  OAI21 U1538 ( .A0(n1120), .A1(n1312), .B0(n1307), .Y(n1309) );
  NOR3B U1539 ( .AN(n1305), .B(n1118), .C(n1125), .Y(n1310) );
  MX2 U1540 ( .A(n1314), .B(n1315), .S0(n1105), .Y(n175) );
  NOR2B U1541 ( .AN(n1316), .B(n1317), .Y(n1314) );
  MX2 U1542 ( .A(n1318), .B(n1319), .S0(n1096), .Y(n174) );
  OAI21 U1543 ( .A0(n1105), .A1(n1312), .B0(n1320), .Y(n1319) );
  INV U1544 ( .A(n1315), .Y(n1320) );
  OAI21 U1545 ( .A0(n1316), .A1(n1312), .B0(n1307), .Y(n1315) );
  NOR3B U1546 ( .AN(n1316), .B(n1104), .C(n1317), .Y(n1318) );
  MX2 U1547 ( .A(n1321), .B(n1322), .S0(n1154), .Y(n173) );
  NOR2B U1548 ( .AN(n1323), .B(n1317), .Y(n1321) );
  MX2 U1549 ( .A(n1324), .B(n1325), .S0(n1123), .Y(n172) );
  OAI21 U1550 ( .A0(n1157), .A1(n1312), .B0(n1326), .Y(n1325) );
  INV U1551 ( .A(n1322), .Y(n1326) );
  OAI21 U1552 ( .A0(n1323), .A1(n1312), .B0(n1307), .Y(n1322) );
  NOR3B U1553 ( .AN(n1323), .B(n1153), .C(n1317), .Y(n1324) );
  MX2 U1554 ( .A(n1327), .B(n1328), .S0(n1116), .Y(n171) );
  INV U1555 ( .A(n1304), .Y(n1328) );
  NOR2B U1556 ( .AN(n1329), .B(n1317), .Y(n1327) );
  INV U1557 ( .A(n1305), .Y(n1317) );
  OAI2BB2 U1558 ( .B0(n1304), .B1(n1112), .A0N(n1305), .A1N(n1330), .Y(n170)
         );
  NOR2B U1559 ( .AN(n1329), .B(n1115), .Y(n1330) );
  NOR2B U1560 ( .AN(n1307), .B(n1312), .Y(n1305) );
  NOR2B U1561 ( .AN(n1307), .B(n1331), .Y(n1304) );
  NOR2 U1562 ( .A(n1329), .B(n1312), .Y(n1331) );
  INV U1563 ( .A(n1332), .Y(n1312) );
  NOR3B U1564 ( .AN(n1323), .B(n1153), .C(n1122), .Y(n1329) );
  NOR3B U1565 ( .AN(n1316), .B(n1104), .C(n1142), .Y(n1323) );
  NOR3 U1566 ( .A(n1118), .B(n1125), .C(n1085), .Y(n1316) );
  MX2 U1567 ( .A(n1271), .B(n1334), .S0(mode), .Y(n1332) );
  INV U1568 ( .A(sync_right), .Y(n1334) );
  INV U1569 ( .A(graphic_lcd_rst), .Y(n1271) );
  NOR2B U1570 ( .AN(n1114), .B(n1335), .Y(n1333) );
  NOR2 U1571 ( .A(n1117), .B(n1336), .Y(n1335) );
  NOR4 U1572 ( .A(n1085), .B(n1104), .C(n1142), .D(n1337), .Y(n1336) );
  OAI211 U1573 ( .A0(n1121), .A1(n1128), .B0(n1157), .C0(n1124), .Y(n1337) );
  INV U1574 ( .A(n1338), .Y(graphic_lcd_di) );
  MX2 U1575 ( .A(n1339), .B(n1340), .S0(n1220), .Y(n1338) );
  XNOR2 U1576 ( .A(mode), .B(graphic_lcd_cs2), .Y(n1220) );
  INV U1577 ( .A(graphic_lcd_cs1), .Y(graphic_lcd_cs2) );
  OR2 U1578 ( .A(refresh), .B(manual_i), .Y(_0_net_) );
endmodule

