
module traffic ( clk, rst_n, nr, ny, ng, sr, sy, sg, wr, wy, wg, er, ey, eg, 
        nsseg1, nsseg2, weseg1, weseg2 );
  output [7:0] nsseg1;
  output [7:0] nsseg2;
  output [7:0] weseg1;
  output [7:0] weseg2;
  input clk, rst_n;
  output nr, ny, ng, sr, sy, sg, wr, wy, wg, er, ey, eg;
  wire   \*Logic1* , ny, wy, N7, N8, N9, N10, N11, N12, N13, N169, N176, er,
         sr, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277;
  wire   [6:0] cnt;
  assign weseg2[7] = \*Logic1* ;
  assign weseg1[7] = \*Logic1* ;
  assign nsseg2[7] = \*Logic1* ;
  assign nsseg1[7] = \*Logic1* ;
  assign nsseg2[1] = ny;
  assign sy = ny;
  assign weseg2[1] = wy;
  assign ey = wy;
  assign nsseg2[3] = nsseg2[4];
  assign nsseg2[0] = nsseg2[4];
  assign weseg2[3] = weseg2[4];
  assign weseg2[0] = weseg2[4];
  assign ng = N169;
  assign sg = N169;
  assign wg = N176;
  assign eg = N176;
  assign wr = er;
  assign nr = sr;

  DFFRHQ \cnt_reg[0]  ( .D(N7), .CK(clk), .RN(n277), .Q(cnt[0]) );
  DFFRHQ \cnt_reg[1]  ( .D(N8), .CK(clk), .RN(n277), .Q(cnt[1]) );
  DFFRHQ \cnt_reg[2]  ( .D(N9), .CK(clk), .RN(n277), .Q(cnt[2]) );
  DFFRHQ \cnt_reg[3]  ( .D(N10), .CK(clk), .RN(n277), .Q(cnt[3]) );
  DFFRHQ \cnt_reg[4]  ( .D(N11), .CK(clk), .RN(n277), .Q(cnt[4]) );
  DFFRHQ \cnt_reg[5]  ( .D(N12), .CK(clk), .RN(n277), .Q(cnt[5]) );
  DFFRHQ \cnt_reg[6]  ( .D(N13), .CK(clk), .RN(n277), .Q(cnt[6]) );
  INV U187 ( .A(n238), .Y(n158) );
  INV U188 ( .A(n158), .Y(n159) );
  LOGIC_1 U189 ( .LOGIC_1_PIN(\*Logic1* ) );
  NAND2 U190 ( .A(n160), .B(weseg2[2]), .Y(weseg2[6]) );
  OR2 U191 ( .A(weseg2[2]), .B(weseg2[4]), .Y(weseg2[5]) );
  OAI21 U192 ( .A0(n161), .A1(weseg2[2]), .B0(n160), .Y(weseg2[4]) );
  AOI211 U193 ( .A0(n162), .A1(n163), .B0(n164), .C0(n165), .Y(n161) );
  INV U194 ( .A(n166), .Y(n163) );
  NAND2B U195 ( .AN(n167), .B(n168), .Y(weseg2[2]) );
  OR3 U196 ( .A(n169), .B(n170), .C(n171), .Y(weseg1[6]) );
  OR3 U197 ( .A(n169), .B(n171), .C(n172), .Y(weseg1[5]) );
  NAND2B U198 ( .AN(weseg1[3]), .B(n173), .Y(weseg1[4]) );
  OR2 U199 ( .A(n169), .B(weseg1[0]), .Y(weseg1[3]) );
  OAI2BB1 U200 ( .A0N(n174), .A1N(n172), .B0(n160), .Y(weseg1[2]) );
  NOR3 U201 ( .A(n164), .B(n165), .C(n175), .Y(n172) );
  MX2 U202 ( .A(n176), .B(n177), .S0(n166), .Y(n175) );
  NAND2 U203 ( .A(n160), .B(n178), .Y(weseg1[1]) );
  INV U204 ( .A(wy), .Y(n160) );
  OR2 U205 ( .A(n179), .B(n171), .Y(weseg1[0]) );
  NOR4B U206 ( .AN(n180), .B(n169), .C(n181), .D(n170), .Y(n171) );
  NOR2B U207 ( .AN(n174), .B(n182), .Y(n170) );
  AOI21 U208 ( .A0(n166), .A1(n183), .B0(n167), .Y(n182) );
  AOI211 U209 ( .A0(n177), .A1(n176), .B0(n164), .C0(n184), .Y(n181) );
  NOR2 U210 ( .A(n177), .B(n176), .Y(n164) );
  INV U211 ( .A(n162), .Y(n176) );
  NOR2B U212 ( .AN(n185), .B(n173), .Y(n169) );
  NOR2B U213 ( .AN(n178), .B(n179), .Y(n180) );
  AOI22 U214 ( .A0(n185), .A1(n174), .B0(n186), .B1(n187), .Y(n178) );
  INV U215 ( .A(n173), .Y(n186) );
  NAND2 U216 ( .A(n168), .B(n188), .Y(n173) );
  XOR2 U217 ( .A(cnt[0]), .B(n189), .Y(n188) );
  NOR3 U218 ( .A(n167), .B(n162), .C(n190), .Y(n185) );
  MX2 U219 ( .A(n166), .B(n191), .S0(n177), .Y(n190) );
  NOR2 U220 ( .A(n166), .B(n191), .Y(n167) );
  NOR2B U221 ( .AN(n187), .B(n192), .Y(n179) );
  INV U222 ( .A(n174), .Y(n192) );
  AOI211 U223 ( .A0(n189), .A1(N7), .B0(n193), .C0(n184), .Y(n174) );
  INV U224 ( .A(n168), .Y(n184) );
  NOR2 U225 ( .A(cnt[6]), .B(n194), .Y(n168) );
  AOI21 U226 ( .A0(n195), .A1(n196), .B0(n197), .Y(n194) );
  NOR2B U227 ( .AN(n183), .B(n166), .Y(n187) );
  AOI2BB1 U228 ( .A0N(cnt[2]), .A1N(n198), .B0(n199), .Y(n166) );
  NOR2 U229 ( .A(n165), .B(n200), .Y(n183) );
  XNOR2 U230 ( .A(n162), .B(n177), .Y(n200) );
  ADDF U231 ( .A(cnt[1]), .B(n189), .CI(n193), .S(n177) );
  XOR2 U232 ( .A(cnt[3]), .B(n199), .Y(n162) );
  INV U233 ( .A(n191), .Y(n165) );
  ADDF U234 ( .A(cnt[4]), .B(n189), .CI(n195), .S(n191) );
  NOR2 U235 ( .A(cnt[3]), .B(n199), .Y(n195) );
  NOR2 U236 ( .A(n201), .B(n202), .Y(n199) );
  INV U237 ( .A(n198), .Y(n202) );
  NOR2B U238 ( .AN(cnt[1]), .B(n203), .Y(n198) );
  NOR2 U239 ( .A(n189), .B(n193), .Y(n203) );
  NOR2 U240 ( .A(n189), .B(N7), .Y(n193) );
  AOI211 U241 ( .A0(n204), .A1(n196), .B0(n205), .C0(ny), .Y(sr) );
  INV U242 ( .A(n206), .Y(n205) );
  NAND2 U243 ( .A(n207), .B(nsseg2[2]), .Y(nsseg2[6]) );
  OR2 U244 ( .A(nsseg2[2]), .B(nsseg2[4]), .Y(nsseg2[5]) );
  OAI21 U245 ( .A0(n208), .A1(nsseg2[2]), .B0(n207), .Y(nsseg2[4]) );
  AOI211 U246 ( .A0(n209), .A1(n210), .B0(n211), .C0(n212), .Y(n208) );
  NAND2B U247 ( .AN(n213), .B(n214), .Y(nsseg2[2]) );
  OR3 U248 ( .A(n215), .B(n216), .C(n217), .Y(nsseg1[6]) );
  OR3 U249 ( .A(n215), .B(n218), .C(n217), .Y(nsseg1[5]) );
  NAND2B U250 ( .AN(nsseg1[3]), .B(n219), .Y(nsseg1[4]) );
  OR2 U251 ( .A(n215), .B(nsseg1[0]), .Y(nsseg1[3]) );
  OAI2BB1 U252 ( .A0N(n218), .A1N(n220), .B0(n207), .Y(nsseg1[2]) );
  NAND2 U253 ( .A(n207), .B(n221), .Y(nsseg1[1]) );
  INV U254 ( .A(ny), .Y(n207) );
  OR2 U255 ( .A(n222), .B(n217), .Y(nsseg1[0]) );
  NOR4BB U256 ( .AN(n223), .BN(n224), .C(n215), .D(n216), .Y(n217) );
  NOR2 U257 ( .A(n225), .B(n226), .Y(n216) );
  AOI22 U258 ( .A0(n213), .A1(n227), .B0(n228), .B1(n229), .Y(n225) );
  NOR2B U259 ( .AN(n230), .B(n219), .Y(n215) );
  OAI21 U260 ( .A0(n231), .A1(n218), .B0(n214), .Y(n224) );
  NOR3B U261 ( .AN(n232), .B(n211), .C(n212), .Y(n218) );
  MX2 U262 ( .A(n233), .B(n210), .S0(n209), .Y(n232) );
  AOI211 U263 ( .A0(n234), .A1(n227), .B0(n209), .C0(n212), .Y(n231) );
  NOR2B U264 ( .AN(n233), .B(n234), .Y(n212) );
  INV U265 ( .A(n233), .Y(n227) );
  NOR2B U266 ( .AN(n221), .B(n222), .Y(n223) );
  AOI22 U267 ( .A0(n230), .A1(n220), .B0(n235), .B1(n236), .Y(n221) );
  INV U268 ( .A(n219), .Y(n235) );
  NAND2 U269 ( .A(n214), .B(n237), .Y(n219) );
  XNOR2 U270 ( .A(cnt[0]), .B(n159), .Y(n237) );
  INV U271 ( .A(n226), .Y(n220) );
  NOR3B U272 ( .AN(n239), .B(n213), .C(n210), .Y(n230) );
  NOR2B U273 ( .AN(n211), .B(n229), .Y(n213) );
  MX2 U274 ( .A(n211), .B(n209), .S0(n233), .Y(n239) );
  INV U275 ( .A(n229), .Y(n209) );
  NOR2B U276 ( .AN(n236), .B(n226), .Y(n222) );
  OAI211 U277 ( .A0(cnt[0]), .A1(n159), .B0(n214), .C0(n240), .Y(n226) );
  INV U278 ( .A(n241), .Y(n240) );
  NOR2 U279 ( .A(cnt[6]), .B(n242), .Y(n214) );
  AOI21 U280 ( .A0(n196), .A1(n243), .B0(n197), .Y(n242) );
  NOR2B U281 ( .AN(n228), .B(n229), .Y(n236) );
  XNOR2 U282 ( .A(cnt[2]), .B(n244), .Y(n229) );
  NOR2 U283 ( .A(n211), .B(n245), .Y(n228) );
  XNOR2 U284 ( .A(n233), .B(n234), .Y(n245) );
  INV U285 ( .A(n210), .Y(n234) );
  ADDF U286 ( .A(n159), .B(n246), .CI(n247), .S(n210) );
  ADDF U287 ( .A(cnt[1]), .B(n159), .CI(n241), .S(n233) );
  NOR2B U288 ( .AN(n243), .B(n248), .Y(n211) );
  XNOR2 U289 ( .A(cnt[4]), .B(n159), .Y(n248) );
  OAI22 U290 ( .A0(n249), .A1(n247), .B0(cnt[3]), .B1(n159), .Y(n243) );
  OR2 U291 ( .A(cnt[2]), .B(n244), .Y(n247) );
  NOR2B U292 ( .AN(cnt[1]), .B(n250), .Y(n244) );
  NOR2B U293 ( .AN(n159), .B(n241), .Y(n250) );
  NOR2B U294 ( .AN(n159), .B(N7), .Y(n241) );
  NOR2B U295 ( .AN(n159), .B(n246), .Y(n249) );
  NOR2B U296 ( .AN(n251), .B(n252), .Y(n238) );
  OAI2BB1 U297 ( .A0N(n253), .A1N(n254), .B0(cnt[4]), .Y(n251) );
  INV U298 ( .A(rst_n), .Y(n277) );
  NOR4B U299 ( .AN(n255), .B(n256), .C(N176), .D(wy), .Y(er) );
  NOR2B U300 ( .AN(n257), .B(cnt[4]), .Y(n256) );
  XNOR2 U301 ( .A(cnt[2]), .B(n254), .Y(N9) );
  XNOR2 U302 ( .A(cnt[1]), .B(N7), .Y(N8) );
  INV U303 ( .A(cnt[0]), .Y(N7) );
  NOR3B U304 ( .AN(n258), .B(cnt[6]), .C(n189), .Y(N176) );
  NOR2B U305 ( .AN(n204), .B(n259), .Y(n189) );
  NOR2B U306 ( .AN(cnt[4]), .B(n260), .Y(n259) );
  NOR2 U307 ( .A(cnt[3]), .B(n261), .Y(n260) );
  AOI2BB1 U308 ( .A0N(cnt[1]), .A1N(cnt[0]), .B0(n201), .Y(n261) );
  OAI31 U309 ( .A0(cnt[0]), .A1(cnt[4]), .A2(cnt[3]), .B0(cnt[5]), .Y(n258) );
  OAI2BB2 U310 ( .B0(cnt[0]), .B1(n206), .A0N(n262), .A1N(n263), .Y(N169) );
  NOR2 U311 ( .A(cnt[4]), .B(n257), .Y(n263) );
  NOR4BB U312 ( .AN(n264), .BN(n204), .C(cnt[0]), .D(cnt[3]), .Y(n257) );
  AOI31 U313 ( .A0(cnt[0]), .A1(cnt[2]), .A2(cnt[3]), .B0(n252), .Y(n262) );
  INV U314 ( .A(n204), .Y(n252) );
  XOR2 U315 ( .A(cnt[6]), .B(n265), .Y(N13) );
  NOR2B U316 ( .AN(n266), .B(n267), .Y(n265) );
  XNOR2 U317 ( .A(n266), .B(n267), .Y(N12) );
  NAND2 U318 ( .A(cnt[4]), .B(n268), .Y(n267) );
  NOR2 U319 ( .A(n269), .B(n197), .Y(n266) );
  OAI31 U320 ( .A0(n201), .A1(n254), .A2(n255), .B0(n270), .Y(wy) );
  INV U321 ( .A(n269), .Y(n270) );
  NAND3B U322 ( .AN(cnt[3]), .B(n271), .C(cnt[5]), .Y(n255) );
  OAI2BB2 U323 ( .B0(n254), .B1(n206), .A0N(n272), .A1N(n273), .Y(ny) );
  NOR4B U324 ( .AN(n204), .B(cnt[1]), .C(cnt[0]), .D(cnt[3]), .Y(n273) );
  NOR2B U325 ( .AN(cnt[4]), .B(n201), .Y(n272) );
  INV U326 ( .A(cnt[2]), .Y(n201) );
  NAND3 U327 ( .A(cnt[4]), .B(n204), .C(n253), .Y(n206) );
  NOR2 U328 ( .A(cnt[2]), .B(cnt[3]), .Y(n253) );
  NOR2 U329 ( .A(cnt[6]), .B(cnt[5]), .Y(n204) );
  XNOR2 U330 ( .A(n268), .B(n196), .Y(N11) );
  INV U331 ( .A(cnt[4]), .Y(n196) );
  NOR2B U332 ( .AN(n274), .B(n275), .Y(n268) );
  XNOR2 U333 ( .A(n274), .B(n275), .Y(N10) );
  NAND2B U334 ( .AN(n254), .B(cnt[2]), .Y(n275) );
  NAND2 U335 ( .A(cnt[1]), .B(cnt[0]), .Y(n254) );
  NOR2 U336 ( .A(n269), .B(n246), .Y(n274) );
  NOR4BB U337 ( .AN(n276), .BN(n264), .C(n197), .D(n246), .Y(n269) );
  INV U338 ( .A(cnt[3]), .Y(n246) );
  INV U339 ( .A(cnt[5]), .Y(n197) );
  NOR2 U340 ( .A(cnt[1]), .B(cnt[2]), .Y(n264) );
  NOR2B U341 ( .AN(n271), .B(cnt[0]), .Y(n276) );
  NOR2 U342 ( .A(cnt[6]), .B(cnt[4]), .Y(n271) );
endmodule

