
module gray (RGB, clk, out_gray);
 input [23:0] RGB;
 input clk;
 output [7:0] out_gray;
  wire \net_Buf-pad-RGB[3]_IN_to_RIGHT_I14_54_0 ;
  wire \net_Buf-pad-RGB[3]_RIGHT_H6C2_to_H6E24_50_0 ;
  wire \net_Buf-pad-RGB[3]_S0_F_B1_to_F14_50_0 ;
  wire \net_Buf-pad-RGB[3]_S0_G_B1_to_G14_50_0 ;
  wire \net_Buf-pad-RGB[19]_IN_to_RIGHT_I327_54_0 ;
  wire \net_Buf-pad-RGB[19]_RIGHT_LLV6_to_RIGHT_LLV08_54_0 ;
  wire \net_Buf-pad-RGB[19]_RIGHT_V6N1_to_RIGHT_V6M15_54_0 ;
  wire \net_Buf-pad-RGB[19]_RIGHT_H6W2_to_H6M25_51_0 ;
  wire \net_Buf-pad-RGB[19]_N16_to_S164_51_0 ;
  wire \net_Buf-pad-RGB[19]_W18_to_E184_50_0 ;
  wire \net_Buf-pad-RGB[19]_S0_F_B2_to_F24_50_0 ;
  wire \net_Buf-pad-RGB[19]_S0_G_B2_to_G24_50_0 ;
  wire \net_Lut-U26_0_Y_to_S0_Y4_50_0 ;
  wire \net_Lut-U26_0_H6W1_to_H6M14_47_0 ;
  wire \net_Lut-U26_0_S9_to_N95_47_0 ;
  wire \net_Lut-U26_0_S0_F_B1_to_F15_47_0 ;
  wire net_VCC_Y_to_S0_Y5_47_0;
  wire net_VCC_S0_F_B2_to_F25_47_0;
  wire \net_Buf-pad-clk_GCLKOUT_to_CLKB_CLKPAD135_28_0 ;
  wire \net_Buf-pad-clk_CLKB_GCLKBUF1_IN_to_IN35_28_0 ;
  wire \net_out_gray_reg[7]_XQ_to_S0_XQ5_11_0 ;
  wire \net_out_gray_reg[7]_H6W6_to_H6E65_5_0 ;
  wire \net_out_gray_reg[7]_V6S6_to_V6N611_5_0 ;
  wire \net_out_gray_reg[7]_H6W10_to_LEFT_H6M1011_2_0 ;
  wire \net_out_gray_reg[7]_LEFT_H6B11_to_H6M1111_3_0 ;
  wire \net_out_gray_reg[7]_N23_to_S2310_3_0 ;
  wire \net_out_gray_reg[7]_W1_to_LEFT_E110_2_0 ;
  wire \net_out_gray_reg[7]_LEFT_O1_to_OUT10_2_0 ;
  wire \net_out_gray_reg[6]_YQ_to_S0_YQ5_11_0 ;
  wire \net_out_gray_reg[6]_H6W8_to_H6E85_5_0 ;
  wire \net_out_gray_reg[6]_V6S8_to_V6N811_5_0 ;
  wire \net_out_gray_reg[6]_H6W6_to_LEFT_H6M611_2_0 ;
  wire \net_out_gray_reg[6]_LEFT_H6B7_to_H6M711_3_0 ;
  wire \net_out_gray_reg[6]_N17_to_S1710_3_0 ;
  wire \net_out_gray_reg[6]_W23_to_LEFT_E2310_2_0 ;
  wire \net_out_gray_reg[6]_LEFT_O2_to_OUT10_2_0 ;
  wire \net_out_gray_reg[5]_XQ_to_S0_XQ5_32_0 ;
  wire \net_out_gray_reg[5]_H6W1_to_H6E15_25_0 ;
  wire \net_out_gray_reg[5]_H6W1_to_H6E15_19_0 ;
  wire \net_out_gray_reg[5]_H6W1_to_H6E15_12_0 ;
  wire \net_out_gray_reg[5]_H6W1_to_H6E15_6_0 ;
  wire \net_out_gray_reg[5]_V6S1_to_V6M18_6_0 ;
  wire \net_out_gray_reg[5]_H6W1_to_LEFT_H6B18_2_0 ;
  wire \net_out_gray_reg[5]_LEFT_O1_to_OUT8_2_0 ;
  wire \net_out_gray_reg[4]_YQ_to_S0_YQ5_32_0 ;
  wire \net_out_gray_reg[4]_LLH6_to_LEFT_LLH105_2_0 ;
  wire \net_out_gray_reg[4]_LEFT_H6B0_to_H6M05_3_0 ;
  wire \net_out_gray_reg[4]_V6S0_to_V6M08_3_0 ;
  wire \net_out_gray_reg[4]_S4_to_N49_3_0 ;
  wire \net_out_gray_reg[4]_W9_to_LEFT_E99_2_0 ;
  wire \net_out_gray_reg[4]_LEFT_O1_to_OUT9_2_0 ;
  wire \net_out_gray_reg[3]_XQ_to_S0_XQ4_11_0 ;
  wire \net_out_gray_reg[3]_LLH6_to_LLH04_5_0 ;
  wire \net_out_gray_reg[3]_H6W1_to_LEFT_H6M14_2_0 ;
  wire \net_out_gray_reg[3]_LEFT_O1_to_OUT4_2_0 ;
  wire \net_out_gray_reg[2]_YQ_to_S0_YQ4_11_0 ;
  wire \net_out_gray_reg[2]_H6W6_to_H6E64_5_0 ;
  wire \net_out_gray_reg[2]_H6W6_to_LEFT_H6M64_2_0 ;
  wire \net_out_gray_reg[2]_LEFT_H6B7_to_H6M74_3_0 ;
  wire \net_out_gray_reg[2]_S16_to_N165_3_0 ;
  wire \net_out_gray_reg[2]_W21_to_LEFT_E215_2_0 ;
  wire \net_out_gray_reg[2]_LEFT_O3_to_OUT5_2_0 ;
  wire \net_out_gray_reg[1]_XQ_to_S0_XQ6_16_0 ;
  wire \net_out_gray_reg[1]_LLH6_to_LLH06_9_0 ;
  wire \net_out_gray_reg[1]_H6W0_to_H6E06_3_0 ;
  wire \net_out_gray_reg[1]_W5_to_LEFT_E56_2_0 ;
  wire \net_out_gray_reg[1]_LEFT_O1_to_OUT6_2_0 ;
  wire \net_out_gray_reg[0]_YQ_to_S0_YQ6_16_0 ;
  wire \net_out_gray_reg[0]_LLH0_to_LLH66_9_0 ;
  wire \net_out_gray_reg[0]_H6W2_to_H6E26_3_0 ;
  wire \net_out_gray_reg[0]_W17_to_LEFT_E176_2_0 ;
  wire \net_out_gray_reg[0]_LEFT_O2_to_OUT6_2_0 ;
  wire net_U3_CO_COUT_to_CO_1_LOCAL3_35_0;
  wire net_U3_CO_LLH6_to_LLH63_9_0;
  wire net_U3_CO_H6E3_to_H6M33_12_0;
  wire net_U3_CO_V6S3_to_V6M36_12_0;
  wire net_U3_CO_W20_to_E206_11_0;
  wire net_U3_CO_N0_to_S05_11_0;
  wire net_U3_CO_S0_BX_B_to_BX5_11_0;
  wire \net_IBuf-clkpad-clk_OUT_to_CLKB_GCLK1_PW35_28_0 ;
  wire \net_IBuf-clkpad-clk_CLKB_GCLK1_to_CLKC_GCLK118_28_0 ;
  wire \net_IBuf-clkpad-clk_CLKC_HGCLK1_to_BRAM_CLKH_GCLK118_1_0 ;
  wire \net_IBuf-clkpad-clk_BRAM_CLKH_VGCLK1_to_BRAM_GCLKIN15_1_0 ;
  wire \net_IBuf-clkpad-clk_BRAM_GCLK_CLBD1_to_GCLK15_11_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK5_11_0 ;
  wire \net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK15_28_0 ;
  wire \net_IBuf-clkpad-clk_CLKV_GCLK_BUFR1_to_GCLK15_32_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK5_32_0 ;
  wire \net_IBuf-clkpad-clk_BRAM_GCLK_CLBC1_to_GCLK14_11_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK4_11_0 ;
  wire \net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK16_16_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK6_16_0 ;
  wire net_U4_S_X_to_S0_X3_35_0;
  wire net_U4_S_LLH0_to_LLH03_9_0;
  wire net_U4_S_H6E0_to_H6M03_12_0;
  wire net_U4_S_V6S0_to_V6M06_12_0;
  wire net_U4_S_W3_to_E36_11_0;
  wire net_U4_S_N3_to_S35_11_0;
  wire net_U4_S_S0_BY_B_to_BY5_11_0;
  wire net_U7_S_Y_to_S1_Y3_40_0;
  wire net_U7_S_H6W2_to_H6E23_34_0;
  wire net_U7_S_H6W2_to_H6M23_31_0;
  wire net_U7_S_V6S2_to_V6M26_31_0;
  wire net_U7_S_E13_to_W136_32_0;
  wire net_U7_S_N8_to_S85_32_0;
  wire net_U7_S_S0_BX_B_to_BX5_32_0;
  wire net_U11_S_Y_to_S1_Y3_42_0;
  wire net_U11_S_H6W4_to_H6E43_35_0;
  wire net_U11_S_H6W4_to_H6M43_32_0;
  wire net_U11_S_S2_to_N24_32_0;
  wire net_U11_S_S2_to_N25_32_0;
  wire net_U11_S_S0_BY_B_to_BY5_32_0;
  wire net_U15_S_Y_to_S1_Y4_42_0;
  wire net_U15_S_LLH0_to_LLH64_9_0;
  wire net_U15_S_H6E3_to_H6M34_12_0;
  wire net_U15_S_W3_to_E34_11_0;
  wire net_U15_S_S0_BX_B_to_BX4_11_0;
  wire net_U19_S_X_to_S0_X4_44_0;
  wire net_U19_S_LLH6_to_LLH04_11_0;
  wire net_U19_S_S0_BY_B_to_BY4_11_0;
  wire net_U24_S_X_to_S1_X5_44_0;
  wire net_U24_S_LLH6_to_LLH65_18_0;
  wire net_U24_S_H6W2_to_H6M25_14_0;
  wire net_U24_S_S18_to_N186_14_0;
  wire net_U24_S_E14_to_W146_16_0;
  wire net_U24_S_S0_BX_B_to_BX6_16_0;
  wire net_U27_S_X_to_S0_X5_45_0;
  wire net_U27_S_LLH0_to_LLH05_19_0;
  wire net_U27_S_H6W0_to_H6M05_16_0;
  wire net_U27_S_S6_to_N66_16_0;
  wire net_U27_S_S0_BY_B_to_BY6_16_0;
  wire \net_Buf-pad-RGB[15]_IN_to_TOP_I11_21_0 ;
  wire \net_Buf-pad-RGB[15]_TOP_H6E2_to_TOP_H6W21_27_0 ;
  wire \net_Buf-pad-RGB[15]_TOP_H6E2_to_TOP_H6W21_34_0 ;
  wire \net_Buf-pad-RGB[15]_TOP_V6D8_to_V6M83_34_0 ;
  wire \net_Buf-pad-RGB[15]_E9_to_W93_35_0 ;
  wire \net_Buf-pad-RGB[15]_S1_G_B1_to_G13_35_0 ;
  wire \net_Buf-pad-RGB[15]_TOP_H6E1_to_TOP_H6W11_27_0 ;
  wire \net_Buf-pad-RGB[15]_TOP_H6E1_to_TOP_H6W11_34_0 ;
  wire \net_Buf-pad-RGB[15]_TOP_V6D10_to_V6M103_34_0 ;
  wire \net_Buf-pad-RGB[15]_E21_to_W213_35_0 ;
  wire \net_Buf-pad-RGB[15]_S0_F_B1_to_F13_35_0 ;
  wire net_U6_CO_COUT_to_CO_0_LOCAL3_42_0;
  wire net_U6_CO_H6W10_to_H6E103_35_0;
  wire net_U6_CO_S1_G_B2_to_G23_35_0;
  wire net_U6_CO_S0_F_B2_to_F23_35_0;
  wire net_U5_CO_XB_to_S1_XB3_35_0;
  wire net_U5_CO_S0_BX_B_to_BX3_35_0;
  wire \net_Buf-pad-RGB[14]_IN_to_TOP_I11_35_0 ;
  wire \net_Buf-pad-RGB[14]_TOP_V6D0_to_V6M03_35_0 ;
  wire \net_Buf-pad-RGB[14]_S1_F_B1_to_F13_35_0 ;
  wire \net_Buf-pad-RGB[14]_TOP_H6E2_to_TOP_H6M21_38_0 ;
  wire \net_Buf-pad-RGB[14]_TOP_V6D10_to_V6M103_38_0 ;
  wire \net_Buf-pad-RGB[14]_E21_to_W213_39_0 ;
  wire \net_Buf-pad-RGB[14]_S0_F_B1_to_F13_39_0 ;
  wire \net_Buf-pad-RGB[7]_IN_to_TOP_I21_48_0 ;
  wire \net_Buf-pad-RGB[7]_TOP_H6W3_to_TOP_H6E31_42_0 ;
  wire \net_Buf-pad-RGB[7]_TOP_H6W3_to_TOP_H6E31_35_0 ;
  wire \net_Buf-pad-RGB[7]_TOP_V6D10_to_V6M103_35_0 ;
  wire \net_Buf-pad-RGB[7]_S1_F_B2_to_F23_35_0 ;
  wire \net_Buf-pad-RGB[7]_TOP_H6W0_to_TOP_H6E01_42_0 ;
  wire \net_Buf-pad-RGB[7]_TOP_H6W0_to_TOP_H6M01_38_0 ;
  wire \net_Buf-pad-RGB[7]_TOP_V6D6_to_V6M63_38_0 ;
  wire \net_Buf-pad-RGB[7]_E12_to_W123_39_0 ;
  wire \net_Buf-pad-RGB[7]_S0_F_B2_to_F23_39_0 ;
  wire \net_Buf-pad-RGB[23]_IN_to_RIGHT_I234_54_0 ;
  wire \net_Buf-pad-RGB[23]_RIGHT_LLV6_to_RIGHT_LLV03_54_0 ;
  wire \net_Buf-pad-RGB[23]_RIGHT_H6W8_to_H6E83_48_0 ;
  wire \net_Buf-pad-RGB[23]_H6W8_to_H6E83_42_0 ;
  wire \net_Buf-pad-RGB[23]_H6W8_to_H6E83_35_0 ;
  wire \net_Buf-pad-RGB[23]_S1_BX_B_to_BX3_35_0 ;
  wire \net_Buf-pad-RGB[23]_RIGHT_H6W4_to_H6E43_48_0 ;
  wire \net_Buf-pad-RGB[23]_H6W4_to_H6E43_42_0 ;
  wire \net_Buf-pad-RGB[23]_W3_to_E33_40_0 ;
  wire \net_Buf-pad-RGB[23]_W3_to_E33_39_0 ;
  wire \net_Buf-pad-RGB[23]_S0_BX_B_to_BX3_39_0 ;
  wire net_U10_S_X_to_S0_X3_39_0;
  wire net_U10_S_E14_to_W143_40_0;
  wire net_U10_S_S1_G_B1_to_G13_40_0;
  wire net_U10_S_E17_to_W173_40_0;
  wire net_U10_S_E17_to_W173_42_0;
  wire net_U10_S_S0_G_B1_to_G13_42_0;
  wire net_U8_CO_XB_to_S1_XB3_40_0;
  wire net_U8_CO_E20_to_W203_42_0;
  wire net_U8_CO_S0_G_B2_to_G23_42_0;
  wire net_U9_CO_XB_to_S0_XB3_42_0;
  wire net_U9_CO_W10_to_E103_40_0;
  wire net_U9_CO_S1_G_B2_to_G23_40_0;
  wire \net_Buf-pad-RGB[13]_IN_to_TOP_I21_40_0 ;
  wire \net_Buf-pad-RGB[13]_TOP_V6B0_to_V6N03_40_0 ;
  wire \net_Buf-pad-RGB[13]_S1_F_B1_to_F13_40_0 ;
  wire \net_Buf-pad-RGB[13]_TOP_V6A3_to_V6N32_40_0 ;
  wire \net_Buf-pad-RGB[13]_S22_to_N223_40_0 ;
  wire \net_Buf-pad-RGB[13]_S0_F_B1_to_F13_40_0 ;
  wire \net_Buf-pad-RGB[6]_IN_to_TOP_I11_50_0 ;
  wire \net_Buf-pad-RGB[6]_TOP_H6W2_to_TOP_H6E21_44_0 ;
  wire \net_Buf-pad-RGB[6]_TOP_H6W2_to_TOP_H6M21_40_0 ;
  wire \net_Buf-pad-RGB[6]_TOP_V6D10_to_V6M103_40_0 ;
  wire \net_Buf-pad-RGB[6]_S1_F_B2_to_F23_40_0 ;
  wire \net_Buf-pad-RGB[6]_TOP_S16_to_N162_40_0 ;
  wire \net_Buf-pad-RGB[6]_S16_to_N163_40_0 ;
  wire \net_Buf-pad-RGB[6]_S0_F_B2_to_F23_40_0 ;
  wire \net_Buf-pad-RGB[22]_IN_to_RIGHT_I330_54_0 ;
  wire \net_Buf-pad-RGB[22]_RIGHT_LLV6_to_RIGHT_LLV65_54_0 ;
  wire \net_Buf-pad-RGB[22]_RIGHT_V6N2_to_RIGHT_V6M22_54_0 ;
  wire \net_Buf-pad-RGB[22]_RIGHT_H6W10_to_H6E102_48_0 ;
  wire \net_Buf-pad-RGB[22]_H6W10_to_H6E102_42_0 ;
  wire \net_Buf-pad-RGB[22]_W23_to_E232_40_0 ;
  wire \net_Buf-pad-RGB[22]_S21_to_N213_40_0 ;
  wire \net_Buf-pad-RGB[22]_S1_BX_B_to_BX3_40_0 ;
  wire \net_Buf-pad-RGB[22]_RIGHT_V6N3_to_RIGHT_V6M32_54_0 ;
  wire \net_Buf-pad-RGB[22]_RIGHT_H6W8_to_H6E82_48_0 ;
  wire \net_Buf-pad-RGB[22]_H6W8_to_H6E82_42_0 ;
  wire \net_Buf-pad-RGB[22]_W11_to_E112_40_0 ;
  wire \net_Buf-pad-RGB[22]_S9_to_N93_40_0 ;
  wire \net_Buf-pad-RGB[22]_S0_BX_B_to_BX3_40_0 ;
  wire net_U14_S_X_to_S0_X3_40_0;
  wire net_U14_S_E11_to_W113_42_0;
  wire net_U14_S_S1_G_B1_to_G13_42_0;
  wire net_U14_S_OUT1_to_OUT_W13_42_0;
  wire net_U14_S_S0_F_B1_to_F13_42_0;
  wire net_U12_CO_XB_to_S1_XB3_42_0;
  wire net_U12_CO_S0_F_B2_to_F23_42_0;
  wire net_U13_CO_COUT_to_CO_0_LOCAL4_42_0;
  wire net_U13_CO_CO_0_to_CIN4_42_0;
  wire \net_Buf-pad-RGB[12]_IN_to_TOP_I11_40_0 ;
  wire \net_Buf-pad-RGB[12]_TOP_V6D0_to_V6M03_40_0 ;
  wire \net_Buf-pad-RGB[12]_E1_to_W13_42_0 ;
  wire \net_Buf-pad-RGB[12]_S1_F_B1_to_F13_42_0 ;
  wire \net_Buf-pad-RGB[12]_TOP_H6E0_to_TOP_H6M01_44_0 ;
  wire \net_Buf-pad-RGB[12]_TOP_V6D6_to_V6M63_44_0 ;
  wire \net_Buf-pad-RGB[12]_W14_to_E143_43_0 ;
  wire \net_Buf-pad-RGB[12]_S0_F_B1_to_F13_43_0 ;
  wire \net_Buf-pad-RGB[5]_IN_to_TOP_I21_53_0 ;
  wire \net_Buf-pad-RGB[5]_TOP_H6W4_to_TOP_H6E41_47_0 ;
  wire \net_Buf-pad-RGB[5]_TOP_H6W4_to_TOP_H6A41_42_0 ;
  wire \net_Buf-pad-RGB[5]_TOP_LLV11_to_LLV02_42_0 ;
  wire \net_Buf-pad-RGB[5]_S2_to_N23_42_0 ;
  wire \net_Buf-pad-RGB[5]_S1_F_B2_to_F23_42_0 ;
  wire \net_Buf-pad-RGB[5]_TOP_H6W3_to_TOP_H6E31_47_0 ;
  wire \net_Buf-pad-RGB[5]_TOP_H6W3_to_TOP_H6M31_44_0 ;
  wire \net_Buf-pad-RGB[5]_TOP_V6D8_to_V6M83_44_0 ;
  wire \net_Buf-pad-RGB[5]_W13_to_E133_43_0 ;
  wire \net_Buf-pad-RGB[5]_S0_F_B2_to_F23_43_0 ;
  wire \net_Buf-pad-RGB[21]_IN_to_RIGHT_I230_54_0 ;
  wire \net_Buf-pad-RGB[21]_RIGHT_LLV0_to_RIGHT_LLV05_54_0 ;
  wire \net_Buf-pad-RGB[21]_RIGHT_V6N0_to_RIGHT_V6M02_54_0 ;
  wire \net_Buf-pad-RGB[21]_RIGHT_H6W6_to_H6E62_48_0 ;
  wire \net_Buf-pad-RGB[21]_H6W6_to_H6E62_42_0 ;
  wire \net_Buf-pad-RGB[21]_S15_to_N153_42_0 ;
  wire \net_Buf-pad-RGB[21]_S1_BX_B_to_BX3_42_0 ;
  wire \net_Buf-pad-RGB[21]_RIGHT_V6N1_to_RIGHT_V6M12_54_0 ;
  wire \net_Buf-pad-RGB[21]_RIGHT_H6D4_to_H6E42_49_0 ;
  wire \net_Buf-pad-RGB[21]_H6W4_to_H6E42_43_0 ;
  wire \net_Buf-pad-RGB[21]_S3_to_N33_43_0 ;
  wire \net_Buf-pad-RGB[21]_S0_BX_B_to_BX3_43_0 ;
  wire net_U18_S_X_to_S0_X3_43_0;
  wire net_U18_S_S7_to_N74_43_0;
  wire net_U18_S_W8_to_E84_42_0;
  wire net_U18_S_S1_G_B1_to_G14_42_0;
  wire net_U18_S_W11_to_E113_42_0;
  wire net_U18_S_S9_to_N94_42_0;
  wire net_U18_S_S0_G_B1_to_G14_42_0;
  wire net_U16_CO_XB_to_S1_XB4_42_0;
  wire net_U16_CO_S0_G_B2_to_G24_42_0;
  wire net_U17_CO_XB_to_S0_XB4_42_0;
  wire net_U17_CO_S1_G_B2_to_G24_42_0;
  wire \net_Buf-pad-RGB[11]_IN_to_TOP_I21_42_0 ;
  wire \net_Buf-pad-RGB[11]_TOP_V6M2_to_V6N24_42_0 ;
  wire \net_Buf-pad-RGB[11]_S1_F_B1_to_F14_42_0 ;
  wire \net_Buf-pad-RGB[11]_TOP_V6S1_to_V6M14_42_0 ;
  wire \net_Buf-pad-RGB[11]_E7_to_W74_43_0 ;
  wire \net_Buf-pad-RGB[11]_S0_F_B1_to_F14_43_0 ;
  wire \net_Buf-pad-RGB[4]_IN_to_TOP_I11_53_0 ;
  wire \net_Buf-pad-RGB[4]_TOP_H6W1_to_TOP_H6E11_47_0 ;
  wire \net_Buf-pad-RGB[4]_TOP_H6W1_to_TOP_H6E11_40_0 ;
  wire \net_Buf-pad-RGB[4]_TOP_V6S6_to_V6M64_40_0 ;
  wire \net_Buf-pad-RGB[4]_E12_to_W124_42_0 ;
  wire \net_Buf-pad-RGB[4]_S1_F_B2_to_F24_42_0 ;
  wire \net_Buf-pad-RGB[4]_TOP_V6S2_to_V6M24_44_0 ;
  wire \net_Buf-pad-RGB[4]_W15_to_E154_43_0 ;
  wire \net_Buf-pad-RGB[4]_S0_F_B2_to_F24_43_0 ;
  wire \net_Buf-pad-RGB[20]_IN_to_RIGHT_I328_54_0 ;
  wire \net_Buf-pad-RGB[20]_RIGHT_LLV6_to_UR_LLV41_54_0 ;
  wire \net_Buf-pad-RGB[20]_UR_V6B1_to_RIGHT_V6N13_54_0 ;
  wire \net_Buf-pad-RGB[20]_RIGHT_H6W6_to_H6E63_48_0 ;
  wire \net_Buf-pad-RGB[20]_H6W6_to_H6E63_42_0 ;
  wire \net_Buf-pad-RGB[20]_S15_to_N154_42_0 ;
  wire \net_Buf-pad-RGB[20]_S1_BX_B_to_BX4_42_0 ;
  wire \net_Buf-pad-RGB[20]_RIGHT_H6D4_to_H6E43_49_0 ;
  wire \net_Buf-pad-RGB[20]_H6W4_to_H6E43_43_0 ;
  wire \net_Buf-pad-RGB[20]_S3_to_N34_43_0 ;
  wire \net_Buf-pad-RGB[20]_S0_BX_B_to_BX4_43_0 ;
  wire net_U23_S_X_to_S0_X4_43_0;
  wire net_U23_S_OUT1_to_OUT_W14_44_0;
  wire net_U23_S_S0_F_B1_to_F14_44_0;
  wire net_U23_S_W10_to_E104_42_0;
  wire net_U23_S_S0_F_B1_to_F14_42_0;
  wire \net_Lut-U21_0_0_X_to_S0_X4_50_0 ;
  wire \net_Lut-U21_0_0_H6W3_to_H6E34_44_0 ;
  wire \net_Lut-U21_0_0_S0_F_B2_to_F24_44_0 ;
  wire \net_Lut-U21_0_0_H6W8_to_H6E84_44_0 ;
  wire \net_Lut-U21_0_0_W11_to_E114_43_0 ;
  wire \net_Lut-U21_0_0_W11_to_E114_42_0 ;
  wire \net_Lut-U21_0_0_S0_F_B2_to_F24_42_0 ;
  wire net_U20_CO_COUT_to_CO_0_LOCAL5_44_0;
  wire net_U20_CO_CO_0_to_CIN5_44_0;
  wire net_U20_CO_H6W1_to_H6M15_40_0;
  wire net_U20_CO_N10_to_S104_40_0;
  wire net_U20_CO_E4_to_W44_42_0;
  wire net_U20_CO_S0_BX_B_to_BX4_42_0;
  wire \net_Buf-pad-RGB[10]_IN_to_TOP_I11_44_0 ;
  wire \net_Buf-pad-RGB[10]_TOP_V6M2_to_V6N24_44_0 ;
  wire \net_Buf-pad-RGB[10]_S14_to_N145_44_0 ;
  wire \net_Buf-pad-RGB[10]_S0_G_B1_to_G15_44_0 ;
  wire \net_Buf-pad-RGB[10]_TOP_V6M1_to_V6N14_44_0 ;
  wire \net_Buf-pad-RGB[10]_S10_to_N105_44_0 ;
  wire \net_Buf-pad-RGB[10]_S1_F_B1_to_F15_44_0 ;
  wire \net_Lut-U26_0InvLut_X_to_S0_X5_47_0 ;
  wire \net_Lut-U26_0InvLut_H6W10_to_H6M105_44_0 ;
  wire \net_Lut-U26_0InvLut_S0_G_B2_to_G25_44_0 ;
  wire \net_Lut-U26_0InvLut_H6W6_to_H6M65_44_0 ;
  wire \net_Lut-U26_0InvLut_S1_F_B2_to_F25_44_0 ;
  wire net_U25_CO_XB_to_S0_XB5_44_0;
  wire net_U25_CO_S1_BX_B_to_BX5_44_0;
  wire \net_Buf-pad-RGB[18]_IN_to_RIGHT_I227_54_0 ;
  wire \net_Buf-pad-RGB[18]_RIGHT_LLV0_to_RIGHT_LLV02_54_0 ;
  wire \net_Buf-pad-RGB[18]_RIGHT_V6S0_to_RIGHT_V6M05_54_0 ;
  wire \net_Buf-pad-RGB[18]_RIGHT_H6D6_to_H6E65_49_0 ;
  wire \net_Buf-pad-RGB[18]_H6W6_to_H6E65_43_0 ;
  wire \net_Buf-pad-RGB[18]_E13_to_W135_44_0 ;
  wire \net_Buf-pad-RGB[18]_S0_F_B1_to_F15_44_0 ;
  wire \net_Buf-pad-RGB[18]_RIGHT_V6N3_to_RIGHT_V6M35_54_0 ;
  wire \net_Buf-pad-RGB[18]_RIGHT_H6W0_to_H6E05_48_0 ;
  wire \net_Buf-pad-RGB[18]_H6W0_to_H6M05_45_0 ;
  wire \net_Buf-pad-RGB[18]_S0_F_B1_to_F15_45_0 ;
  wire \net_Buf-pad-RGB[2]_IN_to_RIGHT_I16_54_0 ;
  wire \net_Buf-pad-RGB[2]_RIGHT_H6C2_to_H6E26_50_0 ;
  wire \net_Buf-pad-RGB[2]_H6W2_to_H6E26_44_0 ;
  wire \net_Buf-pad-RGB[2]_N19_to_S195_44_0 ;
  wire \net_Buf-pad-RGB[2]_S0_F_B2_to_F25_44_0 ;
  wire \net_Buf-pad-RGB[2]_RIGHT_H6W0_to_H6E06_48_0 ;
  wire \net_Buf-pad-RGB[2]_H6W0_to_H6M06_45_0 ;
  wire \net_Buf-pad-RGB[2]_N4_to_S45_45_0 ;
  wire \net_Buf-pad-RGB[2]_S0_F_B2_to_F25_45_0 ;
  wire \net_Buf-pad-RGB[9]_IN_to_TOP_I21_47_0 ;
  wire \net_Buf-pad-RGB[9]_TOP_V6S8_to_V6M84_47_0 ;
  wire \net_Buf-pad-RGB[9]_H6W8_to_H6M84_44_0 ;
  wire \net_Buf-pad-RGB[9]_S11_to_N115_44_0 ;
  wire \net_Buf-pad-RGB[9]_S0_BX_B_to_BX5_44_0 ;
  wire \net_Buf-pad-RGB[9]_TOP_V6C2_to_V6N25_47_0 ;
  wire \net_Buf-pad-RGB[9]_W16_to_E165_46_0 ;
  wire \net_Buf-pad-RGB[9]_W1_to_E15_45_0 ;
  wire \net_Buf-pad-RGB[9]_S0_BX_B_to_BX5_45_0 ;
  wire net_U13_CO_boy_net_YB_to_S0_YB4_42_0;
  wire net_U13_CO_boy_net_N0_to_S03_42_0;
  wire net_U13_CO_boy_net_S1_G_B2_to_G23_42_0;


  defparam iSlice__0___inst.bxmux.CONF = "BX";
  defparam iSlice__0___inst.coutused.CONF = "0";
  defparam iSlice__0___inst.cy0f.CONF = "F1";
  defparam iSlice__0___inst.cy0g.CONF = "G1";
  defparam iSlice__0___inst.cyinit.CONF = "BX";
  defparam iSlice__0___inst.cyself.CONF = "F";
  defparam iSlice__0___inst.cyselg.CONF = "G";
  defparam iSlice__0___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__0___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__0___inst.xbused.CONF = "0";
  defparam iSlice__0___inst.ybmux.CONF = "1";
  defparam iSlice__0___inst.f.INIT = 16'h6;
  defparam iSlice__0___inst.g.INIT = 16'h6;
  SLICE iSlice__0___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(\net_Buf-pad-RGB[23]_S1_BX_B_to_BX3_35_0 ),
    .F1(\net_Buf-pad-RGB[14]_S1_F_B1_to_F13_35_0 ),
    .F2(\net_Buf-pad-RGB[7]_S1_F_B2_to_F23_35_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-RGB[15]_S1_G_B1_to_G13_35_0 ),
    .G2(net_U6_CO_S1_G_B2_to_G23_35_0),
    .G3(),
    .G4(),
    .XQ(),
    .X(),
    .F5(),
    .XB(net_U5_CO_XB_to_S1_XB3_35_0),
    .YQ(),
    .Y(),
    .YB(),
    .COUT(net_U3_CO_COUT_to_CO_1_LOCAL3_35_0)
  );

  defparam iSlice__1___inst.bxmux.CONF = "BX";
  defparam iSlice__1___inst.cyinit.CONF = "BX";
  defparam iSlice__1___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__1___inst.fxmux.CONF = "FXOR";
  defparam iSlice__1___inst.xused.CONF = "0";
  defparam iSlice__1___inst.f.INIT = 16'h6;
  SLICE iSlice__1___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(net_U5_CO_S0_BX_B_to_BX3_35_0),
    .F1(\net_Buf-pad-RGB[15]_S0_F_B1_to_F13_35_0 ),
    .F2(net_U6_CO_S0_F_B2_to_F23_35_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(net_U4_S_X_to_S0_X3_35_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__2___inst.bxmux.CONF = "BX";
  defparam iSlice__2___inst.cy0f.CONF = "F1";
  defparam iSlice__2___inst.cyinit.CONF = "BX";
  defparam iSlice__2___inst.cyself.CONF = "F";
  defparam iSlice__2___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__2___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__2___inst.gymux.CONF = "GXOR";
  defparam iSlice__2___inst.xbused.CONF = "0";
  defparam iSlice__2___inst.ybmux.CONF = "1";
  defparam iSlice__2___inst.yused.CONF = "0";
  defparam iSlice__2___inst.f.INIT = 16'h6;
  defparam iSlice__2___inst.g.INIT = 16'h6;
  SLICE iSlice__2___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(\net_Buf-pad-RGB[22]_S1_BX_B_to_BX3_40_0 ),
    .F1(\net_Buf-pad-RGB[13]_S1_F_B1_to_F13_40_0 ),
    .F2(\net_Buf-pad-RGB[6]_S1_F_B2_to_F23_40_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(net_U10_S_S1_G_B1_to_G13_40_0),
    .G2(net_U9_CO_S1_G_B2_to_G23_40_0),
    .G3(),
    .G4(),
    .XQ(),
    .X(),
    .F5(),
    .XB(net_U8_CO_XB_to_S1_XB3_40_0),
    .YQ(),
    .Y(net_U7_S_Y_to_S1_Y3_40_0),
    .YB(),
    .COUT()
  );

  defparam iSlice__3___inst.bxmux.CONF = "BX";
  defparam iSlice__3___inst.cy0f.CONF = "F1";
  defparam iSlice__3___inst.cyinit.CONF = "BX";
  defparam iSlice__3___inst.cyself.CONF = "F";
  defparam iSlice__3___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__3___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__3___inst.gymux.CONF = "GXOR";
  defparam iSlice__3___inst.xbused.CONF = "0";
  defparam iSlice__3___inst.ybmux.CONF = "1";
  defparam iSlice__3___inst.yused.CONF = "0";
  defparam iSlice__3___inst.f.INIT = 16'h6;
  defparam iSlice__3___inst.g.INIT = 16'h6;
  SLICE iSlice__3___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(\net_Buf-pad-RGB[21]_S1_BX_B_to_BX3_42_0 ),
    .F1(\net_Buf-pad-RGB[12]_S1_F_B1_to_F13_42_0 ),
    .F2(\net_Buf-pad-RGB[5]_S1_F_B2_to_F23_42_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(net_U14_S_S1_G_B1_to_G13_42_0),
    .G2(net_U13_CO_boy_net_S1_G_B2_to_G23_42_0),
    .G3(),
    .G4(),
    .XQ(),
    .X(),
    .F5(),
    .XB(net_U12_CO_XB_to_S1_XB3_42_0),
    .YQ(),
    .Y(net_U11_S_Y_to_S1_Y3_42_0),
    .YB(),
    .COUT()
  );

  defparam iSlice__4___inst.bxmux.CONF = "BX";
  defparam iSlice__4___inst.cy0f.CONF = "F1";
  defparam iSlice__4___inst.cyinit.CONF = "BX";
  defparam iSlice__4___inst.cyself.CONF = "F";
  defparam iSlice__4___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__4___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__4___inst.gymux.CONF = "GXOR";
  defparam iSlice__4___inst.xbused.CONF = "0";
  defparam iSlice__4___inst.ybmux.CONF = "1";
  defparam iSlice__4___inst.yused.CONF = "0";
  defparam iSlice__4___inst.f.INIT = 16'h6;
  defparam iSlice__4___inst.g.INIT = 16'h6;
  SLICE iSlice__4___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(\net_Buf-pad-RGB[20]_S1_BX_B_to_BX4_42_0 ),
    .F1(\net_Buf-pad-RGB[11]_S1_F_B1_to_F14_42_0 ),
    .F2(\net_Buf-pad-RGB[4]_S1_F_B2_to_F24_42_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(net_U18_S_S1_G_B1_to_G14_42_0),
    .G2(net_U17_CO_S1_G_B2_to_G24_42_0),
    .G3(),
    .G4(),
    .XQ(),
    .X(),
    .F5(),
    .XB(net_U16_CO_XB_to_S1_XB4_42_0),
    .YQ(),
    .Y(net_U15_S_Y_to_S1_Y4_42_0),
    .YB(),
    .COUT()
  );

  defparam iSlice__5___inst.bxmux.CONF = "BX";
  defparam iSlice__5___inst.coutused.CONF = "0";
  defparam iSlice__5___inst.cy0f.CONF = "F1";
  defparam iSlice__5___inst.cy0g.CONF = "G1";
  defparam iSlice__5___inst.cyinit.CONF = "BX";
  defparam iSlice__5___inst.cyself.CONF = "F";
  defparam iSlice__5___inst.cyselg.CONF = "G";
  defparam iSlice__5___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__5___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__5___inst.xbused.CONF = "0";
  defparam iSlice__5___inst.ybmux.CONF = "1";
  defparam iSlice__5___inst.f.INIT = 16'h6;
  defparam iSlice__5___inst.g.INIT = 16'h6;
  SLICE iSlice__5___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(\net_Buf-pad-RGB[9]_S0_BX_B_to_BX5_44_0 ),
    .F1(\net_Buf-pad-RGB[18]_S0_F_B1_to_F15_44_0 ),
    .F2(\net_Buf-pad-RGB[2]_S0_F_B2_to_F25_44_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-RGB[10]_S0_G_B1_to_G15_44_0 ),
    .G2(\net_Lut-U26_0InvLut_S0_G_B2_to_G25_44_0 ),
    .G3(),
    .G4(),
    .XQ(),
    .X(),
    .F5(),
    .XB(net_U25_CO_XB_to_S0_XB5_44_0),
    .YQ(),
    .Y(),
    .YB(),
    .COUT(net_U20_CO_COUT_to_CO_0_LOCAL5_44_0)
  );

  defparam iSlice__6___inst.cyinit.CONF = "CIN";
  defparam iSlice__6___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__6___inst.fxmux.CONF = "FXOR";
  defparam iSlice__6___inst.xused.CONF = "0";
  defparam iSlice__6___inst.f.INIT = 16'h6;
  SLICE iSlice__6___inst (
    .CIN(net_U20_CO_CO_0_to_CIN5_44_0),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(net_U23_S_S0_F_B1_to_F14_44_0),
    .F2(\net_Lut-U21_0_0_S0_F_B2_to_F24_44_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(net_U19_S_X_to_S0_X4_44_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__7___inst.bxmux.CONF = "BX";
  defparam iSlice__7___inst.cyinit.CONF = "BX";
  defparam iSlice__7___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__7___inst.fxmux.CONF = "FXOR";
  defparam iSlice__7___inst.xused.CONF = "0";
  defparam iSlice__7___inst.f.INIT = 16'h6;
  SLICE iSlice__7___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(net_U25_CO_S1_BX_B_to_BX5_44_0),
    .F1(\net_Buf-pad-RGB[10]_S1_F_B1_to_F15_44_0 ),
    .F2(\net_Lut-U26_0InvLut_S1_F_B2_to_F25_44_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(net_U24_S_X_to_S1_X5_44_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__8___inst.bxmux.CONF = "BX";
  defparam iSlice__8___inst.cyinit.CONF = "BX";
  defparam iSlice__8___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__8___inst.fxmux.CONF = "FXOR";
  defparam iSlice__8___inst.xused.CONF = "0";
  defparam iSlice__8___inst.f.INIT = 16'h6;
  SLICE iSlice__8___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(\net_Buf-pad-RGB[9]_S0_BX_B_to_BX5_45_0 ),
    .F1(\net_Buf-pad-RGB[18]_S0_F_B1_to_F15_45_0 ),
    .F2(\net_Buf-pad-RGB[2]_S0_F_B2_to_F25_45_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(net_U27_S_X_to_S0_X5_45_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__9___inst.bxmux.CONF = "BX";
  defparam iSlice__9___inst.coutused.CONF = "0";
  defparam iSlice__9___inst.cy0f.CONF = "F1";
  defparam iSlice__9___inst.cy0g.CONF = "G1";
  defparam iSlice__9___inst.cyinit.CONF = "BX";
  defparam iSlice__9___inst.cyself.CONF = "F";
  defparam iSlice__9___inst.cyselg.CONF = "G";
  defparam iSlice__9___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__9___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__9___inst.xbused.CONF = "0";
  defparam iSlice__9___inst.ybmux.CONF = "1";
  defparam iSlice__9___inst.f.INIT = 16'h6;
  defparam iSlice__9___inst.g.INIT = 16'h6;
  SLICE iSlice__9___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(net_U20_CO_S0_BX_B_to_BX4_42_0),
    .F1(net_U23_S_S0_F_B1_to_F14_42_0),
    .F2(\net_Lut-U21_0_0_S0_F_B2_to_F24_42_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(net_U18_S_S0_G_B1_to_G14_42_0),
    .G2(net_U16_CO_S0_G_B2_to_G24_42_0),
    .G3(),
    .G4(),
    .XQ(),
    .X(),
    .F5(),
    .XB(net_U17_CO_XB_to_S0_XB4_42_0),
    .YQ(),
    .Y(),
    .YB(net_U13_CO_boy_net_YB_to_S0_YB4_42_0),
    .COUT(net_U13_CO_COUT_to_CO_0_LOCAL4_42_0)
  );

  defparam iSlice__10___inst.coutused.CONF = "0";
  defparam iSlice__10___inst.cy0f.CONF = "F1";
  defparam iSlice__10___inst.cy0g.CONF = "G1";
  defparam iSlice__10___inst.cyinit.CONF = "CIN";
  defparam iSlice__10___inst.cyself.CONF = "F";
  defparam iSlice__10___inst.cyselg.CONF = "G";
  defparam iSlice__10___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__10___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__10___inst.xbused.CONF = "0";
  defparam iSlice__10___inst.ybmux.CONF = "1";
  defparam iSlice__10___inst.f.INIT = 16'h6;
  defparam iSlice__10___inst.g.INIT = 16'h6;
  SLICE iSlice__10___inst (
    .CIN(net_U13_CO_CO_0_to_CIN4_42_0),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(net_U14_S_S0_F_B1_to_F13_42_0),
    .F2(net_U12_CO_S0_F_B2_to_F23_42_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(net_U10_S_S0_G_B1_to_G13_42_0),
    .G2(net_U8_CO_S0_G_B2_to_G23_42_0),
    .G3(),
    .G4(),
    .XQ(),
    .X(),
    .F5(),
    .XB(net_U9_CO_XB_to_S0_XB3_42_0),
    .YQ(),
    .Y(),
    .YB(),
    .COUT(net_U6_CO_COUT_to_CO_0_LOCAL3_42_0)
  );

  defparam iSlice__11___inst.bxmux.CONF = "BX";
  defparam iSlice__11___inst.cyinit.CONF = "BX";
  defparam iSlice__11___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__11___inst.fxmux.CONF = "FXOR";
  defparam iSlice__11___inst.xused.CONF = "0";
  defparam iSlice__11___inst.f.INIT = 16'h6;
  SLICE iSlice__11___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(\net_Buf-pad-RGB[23]_S0_BX_B_to_BX3_39_0 ),
    .F1(\net_Buf-pad-RGB[14]_S0_F_B1_to_F13_39_0 ),
    .F2(\net_Buf-pad-RGB[7]_S0_F_B2_to_F23_39_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(net_U10_S_X_to_S0_X3_39_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__12___inst.bxmux.CONF = "BX";
  defparam iSlice__12___inst.cyinit.CONF = "BX";
  defparam iSlice__12___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__12___inst.fxmux.CONF = "FXOR";
  defparam iSlice__12___inst.xused.CONF = "0";
  defparam iSlice__12___inst.f.INIT = 16'h6;
  SLICE iSlice__12___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(\net_Buf-pad-RGB[22]_S0_BX_B_to_BX3_40_0 ),
    .F1(\net_Buf-pad-RGB[13]_S0_F_B1_to_F13_40_0 ),
    .F2(\net_Buf-pad-RGB[6]_S0_F_B2_to_F23_40_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(net_U14_S_X_to_S0_X3_40_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__13___inst.bxmux.CONF = "BX";
  defparam iSlice__13___inst.cyinit.CONF = "BX";
  defparam iSlice__13___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__13___inst.fxmux.CONF = "FXOR";
  defparam iSlice__13___inst.xused.CONF = "0";
  defparam iSlice__13___inst.f.INIT = 16'h6;
  SLICE iSlice__13___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(\net_Buf-pad-RGB[21]_S0_BX_B_to_BX3_43_0 ),
    .F1(\net_Buf-pad-RGB[12]_S0_F_B1_to_F13_43_0 ),
    .F2(\net_Buf-pad-RGB[5]_S0_F_B2_to_F23_43_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(net_U18_S_X_to_S0_X3_43_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__14___inst.bxmux.CONF = "BX";
  defparam iSlice__14___inst.cyinit.CONF = "BX";
  defparam iSlice__14___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*A1)";
  defparam iSlice__14___inst.fxmux.CONF = "FXOR";
  defparam iSlice__14___inst.xused.CONF = "0";
  defparam iSlice__14___inst.f.INIT = 16'h6;
  SLICE iSlice__14___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(\net_Buf-pad-RGB[20]_S0_BX_B_to_BX4_43_0 ),
    .F1(\net_Buf-pad-RGB[11]_S0_F_B1_to_F14_43_0 ),
    .F2(\net_Buf-pad-RGB[4]_S0_F_B2_to_F24_43_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(net_U23_S_X_to_S0_X4_43_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__15___inst.bxmux.CONF = "BX";
  defparam iSlice__15___inst.bymux.CONF = "BY";
  defparam iSlice__15___inst.ckinv.CONF = "1";
  defparam iSlice__15___inst.dxmux.CONF = "0";
  defparam iSlice__15___inst.dymux.CONF = "0";
  defparam iSlice__15___inst.ffx.TYPE = "#FF";
  defparam iSlice__15___inst.ffy.TYPE = "#FF";
  defparam iSlice__15___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__15___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__15___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__15___inst.ffy.SYNC_ATTR = "ASYNC";
  SLICE iSlice__15___inst (
    .CIN(),
    .SR(),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK5_11_0 ),
    .CE(),
    .BX(net_U3_CO_S0_BX_B_to_BX5_11_0),
    .F1(),
    .F2(),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(net_U4_S_S0_BY_B_to_BY5_11_0),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(\net_out_gray_reg[7]_XQ_to_S0_XQ5_11_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_out_gray_reg[6]_YQ_to_S0_YQ5_11_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__16___inst.bxmux.CONF = "BX";
  defparam iSlice__16___inst.bymux.CONF = "BY";
  defparam iSlice__16___inst.ckinv.CONF = "1";
  defparam iSlice__16___inst.dxmux.CONF = "0";
  defparam iSlice__16___inst.dymux.CONF = "0";
  defparam iSlice__16___inst.ffx.TYPE = "#FF";
  defparam iSlice__16___inst.ffy.TYPE = "#FF";
  defparam iSlice__16___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__16___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__16___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__16___inst.ffy.SYNC_ATTR = "ASYNC";
  SLICE iSlice__16___inst (
    .CIN(),
    .SR(),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK5_32_0 ),
    .CE(),
    .BX(net_U7_S_S0_BX_B_to_BX5_32_0),
    .F1(),
    .F2(),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(net_U11_S_S0_BY_B_to_BY5_32_0),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(\net_out_gray_reg[5]_XQ_to_S0_XQ5_32_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_out_gray_reg[4]_YQ_to_S0_YQ5_32_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__17___inst.bxmux.CONF = "BX";
  defparam iSlice__17___inst.bymux.CONF = "BY";
  defparam iSlice__17___inst.ckinv.CONF = "1";
  defparam iSlice__17___inst.dxmux.CONF = "0";
  defparam iSlice__17___inst.dymux.CONF = "0";
  defparam iSlice__17___inst.ffx.TYPE = "#FF";
  defparam iSlice__17___inst.ffy.TYPE = "#FF";
  defparam iSlice__17___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__17___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__17___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__17___inst.ffy.SYNC_ATTR = "ASYNC";
  SLICE iSlice__17___inst (
    .CIN(),
    .SR(),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK4_11_0 ),
    .CE(),
    .BX(net_U15_S_S0_BX_B_to_BX4_11_0),
    .F1(),
    .F2(),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(net_U19_S_S0_BY_B_to_BY4_11_0),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(\net_out_gray_reg[3]_XQ_to_S0_XQ4_11_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_out_gray_reg[2]_YQ_to_S0_YQ4_11_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__18___inst.bxmux.CONF = "BX";
  defparam iSlice__18___inst.bymux.CONF = "BY";
  defparam iSlice__18___inst.ckinv.CONF = "1";
  defparam iSlice__18___inst.dxmux.CONF = "0";
  defparam iSlice__18___inst.dymux.CONF = "0";
  defparam iSlice__18___inst.ffx.TYPE = "#FF";
  defparam iSlice__18___inst.ffy.TYPE = "#FF";
  defparam iSlice__18___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__18___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__18___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__18___inst.ffy.SYNC_ATTR = "ASYNC";
  SLICE iSlice__18___inst (
    .CIN(),
    .SR(),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK6_16_0 ),
    .CE(),
    .BX(net_U24_S_S0_BX_B_to_BX6_16_0),
    .F1(),
    .F2(),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(net_U27_S_S0_BY_B_to_BY6_16_0),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(\net_out_gray_reg[1]_XQ_to_S0_XQ6_16_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_out_gray_reg[0]_YQ_to_S0_YQ6_16_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__19___inst.f.CONF = "#LUT:D=(A2*A1)";
  defparam iSlice__19___inst.fxmux.CONF = "F";
  defparam iSlice__19___inst.g.CONF = "#LUT:D=(A2*A1)+(~A2*~A1)";
  defparam iSlice__19___inst.gymux.CONF = "G";
  defparam iSlice__19___inst.xused.CONF = "0";
  defparam iSlice__19___inst.yused.CONF = "0";
  defparam iSlice__19___inst.f.INIT = 16'h8;
  defparam iSlice__19___inst.g.INIT = 16'h9;
  SLICE iSlice__19___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Buf-pad-RGB[3]_S0_F_B1_to_F14_50_0 ),
    .F2(\net_Buf-pad-RGB[19]_S0_F_B2_to_F24_50_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Buf-pad-RGB[3]_S0_G_B1_to_G14_50_0 ),
    .G2(\net_Buf-pad-RGB[19]_S0_G_B2_to_G24_50_0 ),
    .G3(),
    .G4(),
    .XQ(),
    .X(\net_Lut-U21_0_0_X_to_S0_X4_50_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U26_0_Y_to_S0_Y4_50_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__20___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__20___inst.fxmux.CONF = "F";
  defparam iSlice__20___inst.g.CONF = "#LUT:D=1";
  defparam iSlice__20___inst.gymux.CONF = "G";
  defparam iSlice__20___inst.xused.CONF = "0";
  defparam iSlice__20___inst.yused.CONF = "0";
  defparam iSlice__20___inst.f.INIT = 16'h5;
  defparam iSlice__20___inst.g.INIT = 16'hffff;
  SLICE iSlice__20___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U26_0_S0_F_B1_to_F15_47_0 ),
    .F2(net_VCC_S0_F_B2_to_F25_47_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(\net_Lut-U26_0InvLut_X_to_S0_X5_47_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(net_VCC_Y_to_S0_Y5_47_0),
    .YB(),
    .COUT()
  );

  defparam \out_gray[7]_inst .driveattrbox.CONF = "12";
  defparam \out_gray[7]_inst .ioattrbox.CONF = "LVTTL";
  defparam \out_gray[7]_inst .omux.CONF = "O";
  defparam \out_gray[7]_inst .outmux.CONF = "1";
  defparam \out_gray[7]_inst .slew.CONF = "SLOW";
  IOB \out_gray[7]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_out_gray_reg[7]_LEFT_O1_to_OUT10_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(out_gray[7])
  );

  defparam \out_gray[6]_inst .driveattrbox.CONF = "12";
  defparam \out_gray[6]_inst .ioattrbox.CONF = "LVTTL";
  defparam \out_gray[6]_inst .omux.CONF = "O";
  defparam \out_gray[6]_inst .outmux.CONF = "1";
  defparam \out_gray[6]_inst .slew.CONF = "SLOW";
  IOB \out_gray[6]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_out_gray_reg[6]_LEFT_O2_to_OUT10_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(out_gray[6])
  );

  defparam \out_gray[5]_inst .driveattrbox.CONF = "12";
  defparam \out_gray[5]_inst .ioattrbox.CONF = "LVTTL";
  defparam \out_gray[5]_inst .omux.CONF = "O";
  defparam \out_gray[5]_inst .outmux.CONF = "1";
  defparam \out_gray[5]_inst .slew.CONF = "SLOW";
  IOB \out_gray[5]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_out_gray_reg[5]_LEFT_O1_to_OUT8_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(out_gray[5])
  );

  defparam \out_gray[4]_inst .driveattrbox.CONF = "12";
  defparam \out_gray[4]_inst .ioattrbox.CONF = "LVTTL";
  defparam \out_gray[4]_inst .omux.CONF = "O";
  defparam \out_gray[4]_inst .outmux.CONF = "1";
  defparam \out_gray[4]_inst .slew.CONF = "SLOW";
  IOB \out_gray[4]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_out_gray_reg[4]_LEFT_O1_to_OUT9_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(out_gray[4])
  );

  defparam \out_gray[3]_inst .driveattrbox.CONF = "12";
  defparam \out_gray[3]_inst .ioattrbox.CONF = "LVTTL";
  defparam \out_gray[3]_inst .omux.CONF = "O";
  defparam \out_gray[3]_inst .outmux.CONF = "1";
  defparam \out_gray[3]_inst .slew.CONF = "SLOW";
  IOB \out_gray[3]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_out_gray_reg[3]_LEFT_O1_to_OUT4_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(out_gray[3])
  );

  defparam \out_gray[2]_inst .driveattrbox.CONF = "12";
  defparam \out_gray[2]_inst .ioattrbox.CONF = "LVTTL";
  defparam \out_gray[2]_inst .omux.CONF = "O";
  defparam \out_gray[2]_inst .outmux.CONF = "1";
  defparam \out_gray[2]_inst .slew.CONF = "SLOW";
  IOB \out_gray[2]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_out_gray_reg[2]_LEFT_O3_to_OUT5_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(out_gray[2])
  );

  defparam \out_gray[1]_inst .driveattrbox.CONF = "12";
  defparam \out_gray[1]_inst .ioattrbox.CONF = "LVTTL";
  defparam \out_gray[1]_inst .omux.CONF = "O";
  defparam \out_gray[1]_inst .outmux.CONF = "1";
  defparam \out_gray[1]_inst .slew.CONF = "SLOW";
  IOB \out_gray[1]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_out_gray_reg[1]_LEFT_O1_to_OUT6_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(out_gray[1])
  );

  defparam \out_gray[0]_inst .driveattrbox.CONF = "12";
  defparam \out_gray[0]_inst .ioattrbox.CONF = "LVTTL";
  defparam \out_gray[0]_inst .omux.CONF = "O";
  defparam \out_gray[0]_inst .outmux.CONF = "1";
  defparam \out_gray[0]_inst .slew.CONF = "SLOW";
  IOB \out_gray[0]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_out_gray_reg[0]_LEFT_O2_to_OUT6_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(out_gray[0])
  );

  defparam \RGB[23]_inst .imux.CONF = "1";
  defparam \RGB[23]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[23]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[23]_IN_to_RIGHT_I234_54_0 ),
    .IQ(),
    .PAD(RGB[23])
  );

  defparam \RGB[22]_inst .imux.CONF = "1";
  defparam \RGB[22]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[22]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[22]_IN_to_RIGHT_I330_54_0 ),
    .IQ(),
    .PAD(RGB[22])
  );

  defparam \RGB[21]_inst .imux.CONF = "1";
  defparam \RGB[21]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[21]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[21]_IN_to_RIGHT_I230_54_0 ),
    .IQ(),
    .PAD(RGB[21])
  );

  defparam \RGB[20]_inst .imux.CONF = "1";
  defparam \RGB[20]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[20]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[20]_IN_to_RIGHT_I328_54_0 ),
    .IQ(),
    .PAD(RGB[20])
  );

  defparam \RGB[19]_inst .imux.CONF = "1";
  defparam \RGB[19]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[19]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[19]_IN_to_RIGHT_I327_54_0 ),
    .IQ(),
    .PAD(RGB[19])
  );

  defparam \RGB[18]_inst .imux.CONF = "1";
  defparam \RGB[18]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[18]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[18]_IN_to_RIGHT_I227_54_0 ),
    .IQ(),
    .PAD(RGB[18])
  );

  defparam \RGB[15]_inst .imux.CONF = "1";
  defparam \RGB[15]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[15]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[15]_IN_to_TOP_I11_21_0 ),
    .IQ(),
    .PAD(RGB[15])
  );

  defparam \RGB[14]_inst .imux.CONF = "1";
  defparam \RGB[14]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[14]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[14]_IN_to_TOP_I11_35_0 ),
    .IQ(),
    .PAD(RGB[14])
  );

  defparam \RGB[13]_inst .imux.CONF = "1";
  defparam \RGB[13]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[13]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[13]_IN_to_TOP_I21_40_0 ),
    .IQ(),
    .PAD(RGB[13])
  );

  defparam \RGB[12]_inst .imux.CONF = "1";
  defparam \RGB[12]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[12]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[12]_IN_to_TOP_I11_40_0 ),
    .IQ(),
    .PAD(RGB[12])
  );

  defparam \RGB[11]_inst .imux.CONF = "1";
  defparam \RGB[11]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[11]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[11]_IN_to_TOP_I21_42_0 ),
    .IQ(),
    .PAD(RGB[11])
  );

  defparam \RGB[10]_inst .imux.CONF = "1";
  defparam \RGB[10]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[10]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[10]_IN_to_TOP_I11_44_0 ),
    .IQ(),
    .PAD(RGB[10])
  );

  defparam \RGB[9]_inst .imux.CONF = "1";
  defparam \RGB[9]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[9]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[9]_IN_to_TOP_I21_47_0 ),
    .IQ(),
    .PAD(RGB[9])
  );

  defparam \RGB[7]_inst .imux.CONF = "1";
  defparam \RGB[7]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[7]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[7]_IN_to_TOP_I21_48_0 ),
    .IQ(),
    .PAD(RGB[7])
  );

  defparam \RGB[6]_inst .imux.CONF = "1";
  defparam \RGB[6]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[6]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[6]_IN_to_TOP_I11_50_0 ),
    .IQ(),
    .PAD(RGB[6])
  );

  defparam \RGB[5]_inst .imux.CONF = "1";
  defparam \RGB[5]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[5]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[5]_IN_to_TOP_I21_53_0 ),
    .IQ(),
    .PAD(RGB[5])
  );

  defparam \RGB[4]_inst .imux.CONF = "1";
  defparam \RGB[4]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[4]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[4]_IN_to_TOP_I11_53_0 ),
    .IQ(),
    .PAD(RGB[4])
  );

  defparam \RGB[3]_inst .imux.CONF = "1";
  defparam \RGB[3]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[3]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[3]_IN_to_RIGHT_I14_54_0 ),
    .IQ(),
    .PAD(RGB[3])
  );

  defparam \RGB[2]_inst .imux.CONF = "1";
  defparam \RGB[2]_inst .ioattrbox.CONF = "LVTTL";
  IOB \RGB[2]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-RGB[2]_IN_to_RIGHT_I16_54_0 ),
    .IQ(),
    .PAD(RGB[2])
  );

  defparam iGclk_buf__0___inst.cemux.CONF = "1";
  defparam iGclk_buf__0___inst.disable_attr.CONF = "LOW";
  GCLK iGclk_buf__0___inst (
    .CE(),
    .IN(\net_Buf-pad-clk_CLKB_GCLKBUF1_IN_to_IN35_28_0 ),
    .OUT(\net_IBuf-clkpad-clk_OUT_to_CLKB_GCLK1_PW35_28_0 )
  );

  defparam clk_inst.ioattrbox.CONF = "LVTTL";
  GCLKIOB clk_inst (
    .PAD(clk),
    .GCLKOUT(\net_Buf-pad-clk_GCLKOUT_to_CLKB_CLKPAD135_28_0 )
  );

  IOB \RGB[17]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD()
  );

  IOB \RGB[16]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD()
  );

  IOB \RGB[8]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD()
  );

  IOB \RGB[1]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD()
  );

  IOB \RGB[0]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD()
  );

  defparam GSB_RHT_4_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_4_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_4_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_4_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_4_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6c2.CONF = "01110";
  defparam GSB_RHT_4_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_4_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_4_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_4_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_4_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_4_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_4_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_4_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_4_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_4_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_4_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_4_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_4_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(\net_Buf-pad-RGB[3]_RIGHT_H6C2_to_H6E24_50_0 ),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(),
    .RIGHT_LLV6(),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(\net_Buf-pad-RGB[3]_IN_to_RIGHT_I14_54_0 ),
    .RIGHT_I2(),
    .RIGHT_I3(),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_4_50_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_h6w1.CONF = "0010";
  defparam GSB_CNT_4_50_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_h6w3.CONF = "0001";
  defparam GSB_CNT_4_50_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_h6w8.CONF = "000";
  defparam GSB_CNT_4_50_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_50_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_50_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_out7.CONF = "000111";
  defparam GSB_CNT_4_50_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w17.CONF = "01";
  defparam GSB_CNT_4_50_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_out2.CONF = "000111";
  defparam GSB_CNT_4_50_0_inst.sps_out3.CONF = "001011";
  defparam GSB_CNT_4_50_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s0_f_b1.CONF = "100101111";
  defparam GSB_CNT_4_50_0_inst.sps_s0_f_b2.CONF = "011011111";
  defparam GSB_CNT_4_50_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_50_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_50_0_inst.sps_s0_g_b1.CONF = "100010";
  defparam GSB_CNT_4_50_0_inst.sps_s0_g_b2.CONF = "011100";
  defparam GSB_CNT_4_50_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_50_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_50_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_50_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_50_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_50_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_50_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(\net_Buf-pad-RGB[19]_W18_to_E184_50_0 ),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(\net_Buf-pad-RGB[3]_RIGHT_H6C2_to_H6E24_50_0 ),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_Lut-U26_0_H6W1_to_H6M14_47_0 ),
    .H6W2(),
    .H6W3(\net_Lut-U21_0_0_H6W3_to_H6E34_44_0 ),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(\net_Lut-U21_0_0_H6W8_to_H6E84_44_0 ),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-RGB[3]_S0_F_B1_to_F14_50_0 ),
    .S0_F_B2(\net_Buf-pad-RGB[19]_S0_F_B2_to_F24_50_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Buf-pad-RGB[3]_S0_G_B1_to_G14_50_0 ),
    .S0_G_B2(\net_Buf-pad-RGB[19]_S0_G_B2_to_G24_50_0 ),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U21_0_0_X_to_S0_X4_50_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U26_0_Y_to_S0_Y4_50_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_RHT_27_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_27_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_27_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_27_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_27_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_27_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_27_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_27_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_llv0.CONF = "0011011111";
  defparam GSB_RHT_27_54_0_inst.sps_llv6.CONF = "0001111111";
  defparam GSB_RHT_27_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_27_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_27_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_27_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_27_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_27_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_27_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_27_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_27_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_27_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_27_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_27_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_27_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_27_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_27_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_27_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_27_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(\net_Buf-pad-RGB[18]_RIGHT_LLV0_to_RIGHT_LLV02_54_0 ),
    .RIGHT_LLV6(\net_Buf-pad-RGB[19]_RIGHT_LLV6_to_RIGHT_LLV08_54_0 ),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(\net_Buf-pad-RGB[18]_IN_to_RIGHT_I227_54_0 ),
    .RIGHT_I3(\net_Buf-pad-RGB[19]_IN_to_RIGHT_I327_54_0 ),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_RHT_8_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_8_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_8_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_8_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_8_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_8_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_8_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_8_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_8_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_8_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_8_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_8_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_8_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6n1.CONF = "00111011";
  defparam GSB_RHT_8_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6n3.CONF = "00111011";
  defparam GSB_RHT_8_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_8_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_8_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_8_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_8_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(\net_Buf-pad-RGB[19]_RIGHT_V6N1_to_RIGHT_V6M15_54_0 ),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(\net_Buf-pad-RGB[18]_RIGHT_V6N3_to_RIGHT_V6M35_54_0 ),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(\net_Buf-pad-RGB[19]_RIGHT_LLV6_to_RIGHT_LLV08_54_0 ),
    .RIGHT_LLV6(\net_Buf-pad-RGB[18]_RIGHT_LLV0_to_RIGHT_LLV02_54_0 ),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(),
    .RIGHT_I3(),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_RHT_5_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d6.CONF = "110111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w0.CONF = "0101111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w2.CONF = "0101111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_5_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_5_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_5_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_5_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_5_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_5_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_5_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6n0.CONF = "00111011";
  defparam GSB_RHT_5_54_0_inst.sps_v6n1.CONF = "00111011";
  defparam GSB_RHT_5_54_0_inst.sps_v6n2.CONF = "00111011";
  defparam GSB_RHT_5_54_0_inst.sps_v6n3.CONF = "00111011";
  defparam GSB_RHT_5_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_5_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(\net_Buf-pad-RGB[18]_RIGHT_H6D6_to_H6E65_49_0 ),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(\net_Buf-pad-RGB[18]_RIGHT_H6W0_to_H6E05_48_0 ),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(\net_Buf-pad-RGB[19]_RIGHT_H6W2_to_H6M25_51_0 ),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(\net_Buf-pad-RGB[21]_RIGHT_V6N0_to_RIGHT_V6M02_54_0 ),
    .RIGHT_V6N1(\net_Buf-pad-RGB[21]_RIGHT_V6N1_to_RIGHT_V6M12_54_0 ),
    .RIGHT_V6N2(\net_Buf-pad-RGB[22]_RIGHT_V6N2_to_RIGHT_V6M22_54_0 ),
    .RIGHT_V6N3(\net_Buf-pad-RGB[22]_RIGHT_V6N3_to_RIGHT_V6M32_54_0 ),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(\net_Buf-pad-RGB[18]_RIGHT_V6S0_to_RIGHT_V6M05_54_0 ),
    .RIGHT_V6M1(\net_Buf-pad-RGB[19]_RIGHT_V6N1_to_RIGHT_V6M15_54_0 ),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(\net_Buf-pad-RGB[18]_RIGHT_V6N3_to_RIGHT_V6M35_54_0 ),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(\net_Buf-pad-RGB[21]_RIGHT_LLV0_to_RIGHT_LLV05_54_0 ),
    .RIGHT_LLV6(\net_Buf-pad-RGB[22]_RIGHT_LLV6_to_RIGHT_LLV65_54_0 ),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(),
    .RIGHT_I3(),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_5_51_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_51_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_51_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_n16.CONF = "10";
  defparam GSB_CNT_5_51_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_51_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_51_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_51_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_51_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_51_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_51_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(\net_Buf-pad-RGB[19]_N16_to_S164_51_0 ),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(\net_Buf-pad-RGB[19]_RIGHT_H6W2_to_H6M25_51_0 ),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_51_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_51_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_51_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_51_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_51_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_51_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_51_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s16_w18.CONF = "0";
  defparam GSB_CNT_4_51_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_51_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_51_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(\net_Buf-pad-RGB[19]_W18_to_E184_50_0 ),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(\net_Buf-pad-RGB[19]_N16_to_S164_51_0 ),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_47_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_h6w8.CONF = "001";
  defparam GSB_CNT_4_47_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_47_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_47_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_47_0_inst.sps_s9.CONF = "0";
  defparam GSB_CNT_4_47_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_47_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_47_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_47_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_47_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_47_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(\net_Lut-U26_0_S9_to_N95_47_0 ),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(\net_Lut-U26_0_H6W1_to_H6M14_47_0 ),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(\net_Buf-pad-RGB[9]_H6W8_to_H6M84_44_0 ),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(\net_Buf-pad-RGB[9]_TOP_V6S8_to_V6M84_47_0 ),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_47_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_h6w10.CONF = "000";
  defparam GSB_CNT_5_47_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_h6w6.CONF = "000";
  defparam GSB_CNT_5_47_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_47_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_47_0_inst.sps_out6.CONF = "000111";
  defparam GSB_CNT_5_47_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w16.CONF = "01";
  defparam GSB_CNT_5_47_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e11.CONF = "01";
  defparam GSB_CNT_5_47_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_out3.CONF = "001011";
  defparam GSB_CNT_5_47_0_inst.sps_out4.CONF = "000111";
  defparam GSB_CNT_5_47_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0_f_b1.CONF = "011111110";
  defparam GSB_CNT_5_47_0_inst.sps_s0_f_b2.CONF = "001111101";
  defparam GSB_CNT_5_47_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_47_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_47_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_47_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_47_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_47_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_47_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(\net_Lut-U26_0_S9_to_N95_47_0 ),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(\net_Buf-pad-RGB[9]_W16_to_E165_46_0 ),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_Lut-U26_0InvLut_H6W6_to_H6M65_44_0 ),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(\net_Lut-U26_0InvLut_H6W10_to_H6M105_44_0 ),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(\net_Buf-pad-RGB[9]_TOP_V6C2_to_V6N25_47_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U26_0_S0_F_B1_to_F15_47_0 ),
    .S0_F_B2(net_VCC_S0_F_B2_to_F25_47_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U26_0InvLut_X_to_S0_X5_47_0 ),
    .S0_XB(),
    .S0_Y(net_VCC_Y_to_S0_Y5_47_0),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CLKB_35_28_0_inst.sps_h6d0.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6d1.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6d2.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6d3.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh1.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh10.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh4.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh7.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e0.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e1.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e2.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e3.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.spbu_gclk0.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_gclk1.CONF = "0";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e0.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e1.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e2.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e3.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w0.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w1.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w2.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w3.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.sps_ce0.CONF = "1111";
  defparam GSB_CLKB_35_28_0_inst.sps_ce1.CONF = "1111";
  defparam GSB_CLKB_35_28_0_inst.sps_clkfbl.CONF = "010";
  defparam GSB_CLKB_35_28_0_inst.sps_clkfbr.CONF = "010";
  defparam GSB_CLKB_35_28_0_inst.sps_clkinl.CONF = "011";
  defparam GSB_CLKB_35_28_0_inst.sps_clkinr.CONF = "011";
  defparam GSB_CLKB_35_28_0_inst.sps_gclkbuf0_in.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_gclkbuf1_in.CONF = "011111";
  GSB_CLKB GSB_CLKB_35_28_0_inst (
    .CLKB_H6E0(),
    .CLKB_H6E1(),
    .CLKB_H6E2(),
    .CLKB_H6E3(),
    .CLKB_H6A0(),
    .CLKB_H6A1(),
    .CLKB_H6A2(),
    .CLKB_H6A3(),
    .CLKB_H6B0(),
    .CLKB_H6B1(),
    .CLKB_H6B2(),
    .CLKB_H6B3(),
    .CLKB_H6M0(),
    .CLKB_H6M1(),
    .CLKB_H6M2(),
    .CLKB_H6M3(),
    .CLKB_H6C0(),
    .CLKB_H6C1(),
    .CLKB_H6C2(),
    .CLKB_H6C3(),
    .CLKB_H6D0(),
    .CLKB_H6D1(),
    .CLKB_H6D2(),
    .CLKB_H6D3(),
    .CLKB_LLH1(),
    .CLKB_LLH4(),
    .CLKB_LLH7(),
    .CLKB_LLH10(),
    .CLKB_GCLK0(),
    .CLKB_GCLK1(\net_IBuf-clkpad-clk_CLKB_GCLK1_to_CLKC_GCLK118_28_0 ),
    .CLKB_VGCLK0(),
    .CLKB_VGCLK1(),
    .CLKB_VGCLK2(),
    .CLKB_VGCLK3(),
    .CLKB_HGCLK_E0(),
    .CLKB_HGCLK_E1(),
    .CLKB_HGCLK_E2(),
    .CLKB_HGCLK_E3(),
    .CLKB_HGCLK_W0(),
    .CLKB_HGCLK_W1(),
    .CLKB_HGCLK_W2(),
    .CLKB_HGCLK_W3(),
    .CLKB_CLKINL_1(),
    .CLKB_CLKFBL_1(),
    .CLKB_CLKDVL_1(),
    .CLKB_CLK0L_1(),
    .CLKB_CLK90L_1(),
    .CLKB_CLK180L_1(),
    .CLKB_CLK270L_1(),
    .CLKB_CLK2XL_1(),
    .CLKB_CLK2X90L_1(),
    .CLKB_LOCKEDL_1(),
    .CLKB_CLKINR_1(),
    .CLKB_CLKFBR_1(),
    .CLKB_CLKDVR_1(),
    .CLKB_CLK0R_1(),
    .CLKB_CLK90R_1(),
    .CLKB_CLK180R_1(),
    .CLKB_CLK270R_1(),
    .CLKB_CLK2XR_1(),
    .CLKB_CLK2X90R_1(),
    .CLKB_LOCKEDR_1(),
    .CLKB_CLKPAD0(),
    .CLKB_CLKPAD1(\net_Buf-pad-clk_GCLKOUT_to_CLKB_CLKPAD135_28_0 ),
    .CLKB_GCLKBUF0_IN(),
    .CLKB_GCLK0_PW(),
    .CLKB_CE0(),
    .CLKB_GCLKBUF1_IN(\net_Buf-pad-clk_CLKB_GCLKBUF1_IN_to_IN35_28_0 ),
    .CLKB_GCLK1_PW(\net_IBuf-clkpad-clk_OUT_to_CLKB_GCLK1_PW35_28_0 ),
    .CLKB_CE1(),
    .BOT_CLKINL(),
    .BOT_CLKFBL(),
    .BOT_CLKINR(),
    .BOT_CLKFBR(),
    .DLL1_RST_I(),
    .DLL1_RST_O(),
    .DLL0_RST_I(),
    .DLL0_RST_O()
  );

  defparam GSB_CNT_5_11_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_h6w6.CONF = "000";
  defparam GSB_CNT_5_11_0_inst.sps_h6w8.CONF = "000";
  defparam GSB_CNT_5_11_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_11_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_11_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_out2.CONF = "001110";
  defparam GSB_CNT_5_11_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_out4.CONF = "001101";
  defparam GSB_CNT_5_11_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_s0_bx_b.CONF = "101110";
  defparam GSB_CNT_5_11_0_inst.sps_s0_by_b.CONF = "101101";
  defparam GSB_CNT_5_11_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_5_11_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_11_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_11_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_11_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_11_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_11_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_11_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_11_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_11_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s3_e1.CONF = "0";
  defparam GSB_CNT_5_11_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_11_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_11_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(net_U3_CO_N0_to_S05_11_0),
    .S1(),
    .S2(),
    .S3(net_U4_S_N3_to_S35_11_0),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_out_gray_reg[7]_H6W6_to_H6E65_5_0 ),
    .H6W7(),
    .H6W8(\net_out_gray_reg[6]_H6W8_to_H6E85_5_0 ),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBD1_to_GCLK15_11_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(net_U3_CO_S0_BX_B_to_BX5_11_0),
    .S0_BY_B(net_U4_S_S0_BY_B_to_BY5_11_0),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK5_11_0 ),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_out_gray_reg[7]_XQ_to_S0_XQ5_11_0 ),
    .S0_YQ(\net_out_gray_reg[6]_YQ_to_S0_YQ5_11_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s6.CONF = "101";
  defparam GSB_CNT_5_5_0_inst.sps_v6s8.CONF = "101";
  defparam GSB_CNT_5_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_5_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(\net_out_gray_reg[7]_H6W6_to_H6E65_5_0 ),
    .H6E7(),
    .H6E8(\net_out_gray_reg[6]_H6W8_to_H6E85_5_0 ),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(\net_out_gray_reg[7]_V6S6_to_V6N611_5_0 ),
    .V6S7(),
    .V6S8(\net_out_gray_reg[6]_V6S8_to_V6N811_5_0 ),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w10.CONF = "011";
  defparam GSB_CNT_11_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w6.CONF = "011";
  defparam GSB_CNT_11_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_5_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_out_gray_reg[6]_H6W6_to_LEFT_H6M611_2_0 ),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(\net_out_gray_reg[7]_H6W10_to_LEFT_H6M1011_2_0 ),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(\net_out_gray_reg[7]_V6S6_to_V6N611_5_0 ),
    .V6N7(),
    .V6N8(\net_out_gray_reg[6]_V6S8_to_V6N811_5_0 ),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_11_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_11_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_11_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_11_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_11_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_11_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_11_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_11_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_11_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_11_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_11_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_11_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_11_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_11_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_11_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_11_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(\net_out_gray_reg[6]_LEFT_H6B7_to_H6M711_3_0 ),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(\net_out_gray_reg[7]_LEFT_H6B11_to_H6M1111_3_0 ),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(\net_out_gray_reg[6]_H6W6_to_LEFT_H6M611_2_0 ),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(\net_out_gray_reg[7]_H6W10_to_LEFT_H6M1011_2_0 ),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_11_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n17.CONF = "0";
  defparam GSB_CNT_11_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n23.CONF = "0";
  defparam GSB_CNT_11_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(\net_out_gray_reg[6]_N17_to_S1710_3_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(\net_out_gray_reg[7]_N23_to_S2310_3_0 ),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(\net_out_gray_reg[6]_LEFT_H6B7_to_H6M711_3_0 ),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(\net_out_gray_reg[7]_LEFT_H6B11_to_H6M1111_3_0 ),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s17_w23.CONF = "0";
  defparam GSB_CNT_10_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s23_w1.CONF = "0";
  defparam GSB_CNT_10_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(\net_out_gray_reg[7]_W1_to_LEFT_E110_2_0 ),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(\net_out_gray_reg[6]_W23_to_LEFT_E2310_2_0 ),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(\net_out_gray_reg[6]_N17_to_S1710_3_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(\net_out_gray_reg[7]_N23_to_S2310_3_0 ),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_10_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_10_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_10_2_0_inst.sps_o1.CONF = "110101011";
  defparam GSB_LFT_10_2_0_inst.sps_o2.CONF = "110001110";
  defparam GSB_LFT_10_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_10_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_10_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_10_2_0_inst (
    .LEFT_E23(\net_out_gray_reg[6]_W23_to_LEFT_E2310_2_0 ),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(\net_out_gray_reg[7]_W1_to_LEFT_E110_2_0 ),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_out_gray_reg[7]_LEFT_O1_to_OUT10_2_0 ),
    .LEFT_O2(\net_out_gray_reg[6]_LEFT_O2_to_OUT10_2_0 ),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_5_32_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_h6w1.CONF = "0010";
  defparam GSB_CNT_5_32_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_5_32_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_32_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_32_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_out3.CONF = "001101";
  defparam GSB_CNT_5_32_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_out5.CONF = "001110";
  defparam GSB_CNT_5_32_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_s0_bx_b.CONF = "110111";
  defparam GSB_CNT_5_32_0_inst.sps_s0_by_b.CONF = "101011";
  defparam GSB_CNT_5_32_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_5_32_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_32_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_32_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_32_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_32_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_32_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_32_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_32_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_32_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_32_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_32_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(net_U11_S_S2_to_N25_32_0),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(net_U7_S_N8_to_S85_32_0),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_out_gray_reg[5]_H6W1_to_H6E15_25_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(\net_out_gray_reg[4]_LLH6_to_LEFT_LLH105_2_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFR1_to_GCLK15_32_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(net_U7_S_S0_BX_B_to_BX5_32_0),
    .S0_BY_B(net_U11_S_S0_BY_B_to_BY5_32_0),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK5_32_0 ),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_out_gray_reg[5]_XQ_to_S0_XQ5_32_0 ),
    .S0_YQ(\net_out_gray_reg[4]_YQ_to_S0_YQ5_32_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_25_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_h6w1.CONF = "0000";
  defparam GSB_CNT_5_25_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_25_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_25_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_25_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_25_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_25_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_25_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_25_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_25_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(\net_out_gray_reg[5]_H6W1_to_H6E15_25_0 ),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_out_gray_reg[5]_H6W1_to_H6E15_19_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_19_0_inst.sps_h6w0.CONF = "0001";
  defparam GSB_CNT_5_19_0_inst.sps_h6w1.CONF = "0000";
  defparam GSB_CNT_5_19_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_19_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_19_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_19_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_19_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_19_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_19_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_19_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_19_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(\net_out_gray_reg[5]_H6W1_to_H6E15_19_0 ),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(net_U27_S_H6W0_to_H6M05_16_0),
    .H6W1(\net_out_gray_reg[5]_H6W1_to_H6E15_12_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(net_U27_S_LLH0_to_LLH05_19_0),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_12_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_h6w1.CONF = "0000";
  defparam GSB_CNT_5_12_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_12_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_12_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_12_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_12_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_12_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_12_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_12_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_12_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(\net_out_gray_reg[5]_H6W1_to_H6E15_12_0 ),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_out_gray_reg[5]_H6W1_to_H6E15_6_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_6_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w1.CONF = "0000";
  defparam GSB_CNT_5_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_6_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s1.CONF = "0010";
  defparam GSB_CNT_5_6_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_6_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(\net_out_gray_reg[5]_H6W1_to_H6E15_6_0 ),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(\net_out_gray_reg[5]_V6S1_to_V6M18_6_0 ),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_6_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w1.CONF = "0011";
  defparam GSB_CNT_8_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_6_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_6_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_out_gray_reg[5]_H6W1_to_LEFT_H6B18_2_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_out_gray_reg[5]_V6S1_to_V6M18_6_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_8_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_8_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_8_2_0_inst.sps_o1.CONF = "110111011";
  defparam GSB_LFT_8_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_8_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_8_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_8_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_8_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(\net_out_gray_reg[5]_H6W1_to_LEFT_H6B18_2_0 ),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_out_gray_reg[5]_LEFT_O1_to_OUT8_2_0 ),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_LFT_5_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b0.CONF = "00111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_5_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_5_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_5_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_5_2_0_inst.sps_o3.CONF = "110001011";
  defparam GSB_LFT_5_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_5_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_5_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(\net_out_gray_reg[2]_W21_to_LEFT_E215_2_0 ),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(\net_out_gray_reg[4]_LEFT_H6B0_to_H6M05_3_0 ),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(\net_out_gray_reg[4]_LLH6_to_LEFT_LLH105_2_0 ),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(),
    .LEFT_O3(\net_out_gray_reg[2]_LEFT_O3_to_OUT5_2_0 ),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_5_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s0.CONF = "0011";
  defparam GSB_CNT_5_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n16_w21.CONF = "0";
  defparam GSB_CNT_5_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(\net_out_gray_reg[2]_S16_to_N165_3_0 ),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(\net_out_gray_reg[2]_W21_to_LEFT_E215_2_0 ),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(\net_out_gray_reg[4]_LEFT_H6B0_to_H6M05_3_0 ),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(\net_out_gray_reg[4]_V6S0_to_V6M08_3_0 ),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_h6e0.CONF = "0010";
  defparam GSB_CNT_8_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s4.CONF = "01";
  defparam GSB_CNT_8_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(\net_out_gray_reg[4]_S4_to_N49_3_0 ),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(\net_out_gray_reg[4]_V6S0_to_V6M08_3_0 ),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n4_w9.CONF = "0";
  defparam GSB_CNT_9_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(\net_out_gray_reg[4]_S4_to_N49_3_0 ),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(\net_out_gray_reg[4]_W9_to_LEFT_E99_2_0 ),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_9_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_9_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_9_2_0_inst.sps_o1.CONF = "110001011";
  defparam GSB_LFT_9_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_9_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_9_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_9_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_9_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(\net_out_gray_reg[4]_W9_to_LEFT_E99_2_0 ),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_out_gray_reg[4]_LEFT_O1_to_OUT9_2_0 ),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_4_11_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_h6w6.CONF = "000";
  defparam GSB_CNT_4_11_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_4_11_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_11_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_11_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_h6e1.CONF = "0000";
  defparam GSB_CNT_4_11_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_n6.CONF = "01";
  defparam GSB_CNT_4_11_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_out4.CONF = "001110";
  defparam GSB_CNT_4_11_0_inst.sps_out5.CONF = "001101";
  defparam GSB_CNT_4_11_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_s0_bx_b.CONF = "011101";
  defparam GSB_CNT_4_11_0_inst.sps_s0_by_b.CONF = "110111";
  defparam GSB_CNT_4_11_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_4_11_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_11_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_11_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_11_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_11_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_11_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_11_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_11_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_11_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_11_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_11_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(net_U15_S_W3_to_E34_11_0),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_out_gray_reg[2]_H6W6_to_H6E64_5_0 ),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(net_U19_S_LLH6_to_LLH04_11_0),
    .LLH6(\net_out_gray_reg[3]_LLH6_to_LLH04_5_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBC1_to_GCLK14_11_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(net_U15_S_S0_BX_B_to_BX4_11_0),
    .S0_BY_B(net_U19_S_S0_BY_B_to_BY4_11_0),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK4_11_0 ),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_out_gray_reg[3]_XQ_to_S0_XQ4_11_0 ),
    .S0_YQ(\net_out_gray_reg[2]_YQ_to_S0_YQ4_11_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_h6w1.CONF = "0001";
  defparam GSB_CNT_4_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_h6w6.CONF = "101";
  defparam GSB_CNT_4_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_5_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(\net_out_gray_reg[2]_H6W6_to_H6E64_5_0 ),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_out_gray_reg[3]_H6W1_to_LEFT_H6M14_2_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_out_gray_reg[2]_H6W6_to_LEFT_H6M64_2_0 ),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_out_gray_reg[3]_LLH6_to_LLH04_5_0 ),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_4_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_4_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_4_2_0_inst.sps_o1.CONF = "110110111";
  defparam GSB_LFT_4_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_4_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_4_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_4_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_4_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(\net_out_gray_reg[2]_LEFT_H6B7_to_H6M74_3_0 ),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(\net_out_gray_reg[3]_H6W1_to_LEFT_H6M14_2_0 ),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(\net_out_gray_reg[2]_H6W6_to_LEFT_H6M64_2_0 ),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_out_gray_reg[3]_LEFT_O1_to_OUT4_2_0 ),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_4_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s16.CONF = "10";
  defparam GSB_CNT_4_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(\net_out_gray_reg[2]_S16_to_N165_3_0 ),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(\net_out_gray_reg[2]_LEFT_H6B7_to_H6M74_3_0 ),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_16_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_llh0.CONF = "01";
  defparam GSB_CNT_6_16_0_inst.sps_llh6.CONF = "00";
  defparam GSB_CNT_6_16_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_16_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_16_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_out3.CONF = "001110";
  defparam GSB_CNT_6_16_0_inst.sps_out4.CONF = "001101";
  defparam GSB_CNT_6_16_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_s0_bx_b.CONF = "101101";
  defparam GSB_CNT_6_16_0_inst.sps_s0_by_b.CONF = "110111";
  defparam GSB_CNT_6_16_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_6_16_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_16_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_16_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_16_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_16_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_16_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_16_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_16_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_16_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_16_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_16_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(net_U27_S_S6_to_N66_16_0),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(net_U24_S_E14_to_W146_16_0),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_out_gray_reg[0]_LLH0_to_LLH66_9_0 ),
    .LLH6(\net_out_gray_reg[1]_LLH6_to_LLH06_9_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK16_16_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(net_U24_S_S0_BX_B_to_BX6_16_0),
    .S0_BY_B(net_U27_S_S0_BY_B_to_BY6_16_0),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK6_16_0 ),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_out_gray_reg[1]_XQ_to_S0_XQ6_16_0 ),
    .S0_YQ(\net_out_gray_reg[0]_YQ_to_S0_YQ6_16_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_9_0_inst.sps_h6w0.CONF = "0001";
  defparam GSB_CNT_6_9_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w2.CONF = "0001";
  defparam GSB_CNT_6_9_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_9_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_9_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_9_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(\net_out_gray_reg[1]_H6W0_to_H6E06_3_0 ),
    .H6W1(),
    .H6W2(\net_out_gray_reg[0]_H6W2_to_H6E26_3_0 ),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_out_gray_reg[1]_LLH6_to_LLH06_9_0 ),
    .LLH6(\net_out_gray_reg[0]_LLH0_to_LLH66_9_0 ),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w17.CONF = "01";
  defparam GSB_CNT_6_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w5.CONF = "01";
  defparam GSB_CNT_6_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(\net_out_gray_reg[1]_W5_to_LEFT_E56_2_0 ),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(\net_out_gray_reg[0]_W17_to_LEFT_E176_2_0 ),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(\net_out_gray_reg[1]_H6W0_to_H6E06_3_0 ),
    .H6E1(),
    .H6E2(\net_out_gray_reg[0]_H6W2_to_H6E26_3_0 ),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_6_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_6_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_6_2_0_inst.sps_o1.CONF = "110011011";
  defparam GSB_LFT_6_2_0_inst.sps_o2.CONF = "110011011";
  defparam GSB_LFT_6_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_6_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_6_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_6_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(\net_out_gray_reg[0]_W17_to_LEFT_E176_2_0 ),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(\net_out_gray_reg[1]_W5_to_LEFT_E56_2_0 ),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_out_gray_reg[1]_LEFT_O1_to_OUT6_2_0 ),
    .LEFT_O2(\net_out_gray_reg[0]_LEFT_O2_to_OUT6_2_0 ),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_3_35_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_h6w4.CONF = "101";
  defparam GSB_CNT_3_35_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_llh0.CONF = "01";
  defparam GSB_CNT_3_35_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_3_35_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_35_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_35_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w23.CONF = "01";
  defparam GSB_CNT_3_35_0_inst.sps_w3.CONF = "01";
  defparam GSB_CNT_3_35_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_e21.CONF = "01";
  defparam GSB_CNT_3_35_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n21.CONF = "01";
  defparam GSB_CNT_3_35_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_n6.CONF = "10";
  defparam GSB_CNT_3_35_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_n9.CONF = "01";
  defparam GSB_CNT_3_35_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_out2.CONF = "101101";
  defparam GSB_CNT_3_35_0_inst.sps_out3.CONF = "000111";
  defparam GSB_CNT_3_35_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_out5.CONF = "101110";
  defparam GSB_CNT_3_35_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_s0_bx_b.CONF = "100111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_f_b1.CONF = "010101111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_f_b2.CONF = "011110111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_s1_bx_b.CONF = "101101";
  defparam GSB_CNT_3_35_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s1_f_b1.CONF = "010011111";
  defparam GSB_CNT_3_35_0_inst.sps_s1_f_b2.CONF = "001111101";
  defparam GSB_CNT_3_35_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_35_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_35_0_inst.sps_s1_g_b1.CONF = "100000";
  defparam GSB_CNT_3_35_0_inst.sps_s1_g_b2.CONF = "001000";
  defparam GSB_CNT_3_35_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_35_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_35_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_35_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_35_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_35_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_35_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(\net_Buf-pad-RGB[15]_E9_to_W93_35_0 ),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(\net_Buf-pad-RGB[15]_E21_to_W213_35_0 ),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(net_U11_S_H6W4_to_H6E43_35_0),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(\net_Buf-pad-RGB[23]_H6W8_to_H6E83_35_0 ),
    .H6E9(),
    .H6E10(net_U6_CO_H6W10_to_H6E103_35_0),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(net_U11_S_H6W4_to_H6M43_32_0),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(net_U4_S_LLH0_to_LLH03_9_0),
    .LLH6(net_U3_CO_LLH6_to_LLH63_9_0),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(\net_Buf-pad-RGB[14]_TOP_V6D0_to_V6M03_35_0 ),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(\net_Buf-pad-RGB[7]_TOP_V6D10_to_V6M103_35_0 ),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-RGB[15]_S0_F_B1_to_F13_35_0 ),
    .S0_F_B2(net_U6_CO_S0_F_B2_to_F23_35_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(net_U5_CO_S0_BX_B_to_BX3_35_0),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(net_U4_S_X_to_S0_X3_35_0),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Buf-pad-RGB[14]_S1_F_B1_to_F13_35_0 ),
    .S1_F_B2(\net_Buf-pad-RGB[7]_S1_F_B2_to_F23_35_0 ),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(\net_Buf-pad-RGB[15]_S1_G_B1_to_G13_35_0 ),
    .S1_G_B2(net_U6_CO_S1_G_B2_to_G23_35_0),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(\net_Buf-pad-RGB[23]_S1_BX_B_to_BX3_35_0 ),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(net_U5_CO_XB_to_S1_XB3_35_0),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(net_U3_CO_COUT_to_CO_1_LOCAL3_35_0),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_3_9_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_9_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_9_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_h6e0.CONF = "0000";
  defparam GSB_CNT_3_9_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_h6e3.CONF = "0001";
  defparam GSB_CNT_3_9_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_9_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_9_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_9_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_9_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_9_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_9_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(net_U4_S_H6E0_to_H6M03_12_0),
    .H6E1(),
    .H6E2(),
    .H6E3(net_U3_CO_H6E3_to_H6M33_12_0),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(net_U4_S_LLH0_to_LLH03_9_0),
    .LLH6(net_U3_CO_LLH6_to_LLH63_9_0),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_3_12_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_12_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_12_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_v6s0.CONF = "0011";
  defparam GSB_CNT_3_12_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_v6s3.CONF = "0011";
  defparam GSB_CNT_3_12_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_12_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_12_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_12_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_12_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_12_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_12_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(net_U4_S_H6E0_to_H6M03_12_0),
    .H6M1(),
    .H6M2(),
    .H6M3(net_U3_CO_H6E3_to_H6M33_12_0),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(net_U4_S_V6S0_to_V6M06_12_0),
    .V6S1(),
    .V6S2(),
    .V6S3(net_U3_CO_V6S3_to_V6M36_12_0),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_12_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_12_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_12_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_w20.CONF = "01";
  defparam GSB_CNT_6_12_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w3.CONF = "01";
  defparam GSB_CNT_6_12_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_12_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_12_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_12_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_12_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_12_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_12_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(net_U4_S_W3_to_E36_11_0),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(net_U3_CO_W20_to_E206_11_0),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(net_U4_S_V6S0_to_V6M06_12_0),
    .V6M1(),
    .V6M2(),
    .V6M3(net_U3_CO_V6S3_to_V6M36_12_0),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_11_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_11_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_11_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n0_e20.CONF = "0";
  defparam GSB_CNT_6_11_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n3_e3.CONF = "0";
  defparam GSB_CNT_6_11_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_11_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(net_U4_S_W3_to_E36_11_0),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(net_U3_CO_W20_to_E206_11_0),
    .E21(),
    .E22(),
    .E23(),
    .N0(net_U3_CO_N0_to_S05_11_0),
    .N1(),
    .N2(),
    .N3(net_U4_S_N3_to_S35_11_0),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  GSB_CLKC GSB_CLKC_18_28_0_inst (
    .CLKC_GCLK0(),
    .CLKC_GCLK1(\net_IBuf-clkpad-clk_CLKB_GCLK1_to_CLKC_GCLK118_28_0 ),
    .CLKC_GCLK2(),
    .CLKC_GCLK3(),
    .CLKC_HGCLK0(),
    .CLKC_HGCLK1(\net_IBuf-clkpad-clk_CLKC_HGCLK1_to_BRAM_CLKH_GCLK118_1_0 ),
    .CLKC_HGCLK2(),
    .CLKC_HGCLK3(),
    .CLKC_VGCLK0(),
    .CLKC_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK15_28_0 ),
    .CLKC_VGCLK2(),
    .CLKC_VGCLK3()
  );

  GSB_CLKL GSB_CLKL_18_1_0_inst (
    .BRAM_CLKH_GCLK0(),
    .BRAM_CLKH_GCLK1(\net_IBuf-clkpad-clk_CLKC_HGCLK1_to_BRAM_CLKH_GCLK118_1_0 ),
    .BRAM_CLKH_GCLK2(),
    .BRAM_CLKH_GCLK3(),
    .BRAM_CLKH_VGCLK0(),
    .BRAM_CLKH_VGCLK1(\net_IBuf-clkpad-clk_BRAM_CLKH_VGCLK1_to_BRAM_GCLKIN15_1_0 ),
    .BRAM_CLKH_VGCLK2(),
    .BRAM_CLKH_VGCLK3()
  );

  defparam GSB_LBRAMD_5_1_0_inst.sps_llv0.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.spbu_gclk_clbd0.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.spbu_gclk_clbd1.CONF = "0";
  defparam GSB_LBRAMD_5_1_0_inst.spbu_gclk_clbd2.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.spbu_gclk_clbd3.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.spbu_gclk_iobd0.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.spbu_gclk_iobd1.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.spbu_gclk_iobd2.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.spbu_gclk_iobd3.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.sps_addra10.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_addra11.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_addra8.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_addra9.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_addrb10.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_addrb11.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_addrb8.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_addrb9.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_dia14.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_dia15.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_dia6.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_dia7.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_dib14.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_dib15.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_dib6.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_dib7.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed0.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed1.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed10.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed11.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed12.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed13.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed14.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed15.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed16.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed17.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed18.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed19.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed2.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed20.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed21.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed22.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed23.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed3.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed4.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed5.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed6.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed7.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed8.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_ed9.CONF = "11";
  defparam GSB_LBRAMD_5_1_0_inst.sps_h6bd0.CONF = "111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_h6bd1.CONF = "111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_h6bd2.CONF = "111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_h6bd3.CONF = "111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_h6md0.CONF = "111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_h6md1.CONF = "111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_h6md2.CONF = "111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_h6md3.CONF = "111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_lhd0.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_lhd3.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_lhd6.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_lhd9.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_llv4.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_llv8.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_raddrs0.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_raddrs12.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_raddrs16.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_raddrs20.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_raddrs24.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_raddrs28.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_raddrs4.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_raddrs8.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_rdins0.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_rdins12.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_rdins16.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_rdins20.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_rdins24.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_rdins28.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_rdins4.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.sps_rdins8.CONF = "111111";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa11_rdouts19.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa11_rdouts2.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa15_rdouts25.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa15_rdouts8.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa3_rdouts1.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa3_rdouts19.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa3_rdouts2.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa3_rdouts20.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa7_rdouts25.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa7_rdouts26.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa7_rdouts7.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_doa7_rdouts8.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob11_rdouts20.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob11_rdouts3.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob15_rdouts26.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob15_rdouts9.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob3_rdouts2.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob3_rdouts20.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob3_rdouts21.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob3_rdouts3.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob7_rdouts26.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob7_rdouts27.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob7_rdouts8.CONF = "1";
  defparam GSB_LBRAMD_5_1_0_inst.tribuf_dob7_rdouts9.CONF = "1";
  GSB_LBRAMD GSB_LBRAMD_5_1_0_inst (
    .BRAM_ED0(),
    .BRAM_ED1(),
    .BRAM_ED2(),
    .BRAM_ED3(),
    .BRAM_ED4(),
    .BRAM_ED5(),
    .BRAM_ED6(),
    .BRAM_ED7(),
    .BRAM_ED8(),
    .BRAM_ED9(),
    .BRAM_ED10(),
    .BRAM_ED11(),
    .BRAM_ED12(),
    .BRAM_ED13(),
    .BRAM_ED14(),
    .BRAM_ED15(),
    .BRAM_ED16(),
    .BRAM_ED17(),
    .BRAM_ED18(),
    .BRAM_ED19(),
    .BRAM_ED20(),
    .BRAM_ED21(),
    .BRAM_ED22(),
    .BRAM_ED23(),
    .BRAM_H6ED0(),
    .BRAM_H6ED1(),
    .BRAM_H6ED2(),
    .BRAM_H6ED3(),
    .BRAM_H6BD0(),
    .BRAM_H6BD1(),
    .BRAM_H6BD2(),
    .BRAM_H6BD3(),
    .BRAM_H6MD0(),
    .BRAM_H6MD1(),
    .BRAM_H6MD2(),
    .BRAM_H6MD3(),
    .BRAM_H6DD0(),
    .BRAM_H6DD1(),
    .BRAM_H6DD2(),
    .BRAM_H6DD3(),
    .BRAM_LHD0(),
    .BRAM_LHD3(),
    .BRAM_LHD6(),
    .BRAM_LHD9(),
    .BRAM_LLV0(),
    .BRAM_LLV4(),
    .BRAM_LLV8(),
    .BRAM_RDOUTS0(),
    .BRAM_RDOUTS1(),
    .BRAM_RDOUTS2(),
    .BRAM_RDOUTS3(),
    .BRAM_RDOUTS4(),
    .BRAM_RDOUTS7(),
    .BRAM_RDOUTS8(),
    .BRAM_RDOUTS9(),
    .BRAM_RDOUTS12(),
    .BRAM_RDOUTS16(),
    .BRAM_RDOUTS19(),
    .BRAM_RDOUTS20(),
    .BRAM_RDOUTS21(),
    .BRAM_RDOUTS24(),
    .BRAM_RDOUTS25(),
    .BRAM_RDOUTS26(),
    .BRAM_RDOUTS27(),
    .BRAM_RDOUTS28(),
    .BRAM_RADDRS0(),
    .BRAM_RADDRS4(),
    .BRAM_RADDRS8(),
    .BRAM_RADDRS12(),
    .BRAM_RADDRS16(),
    .BRAM_RADDRS17(),
    .BRAM_RADDRS18(),
    .BRAM_RADDRS19(),
    .BRAM_RADDRS20(),
    .BRAM_RADDRS21(),
    .BRAM_RADDRS22(),
    .BRAM_RADDRS23(),
    .BRAM_RADDRS24(),
    .BRAM_RADDRS25(),
    .BRAM_RADDRS26(),
    .BRAM_RADDRS27(),
    .BRAM_RADDRS28(),
    .BRAM_RDINS0(),
    .BRAM_RDINS4(),
    .BRAM_RDINS8(),
    .BRAM_RDINS9(),
    .BRAM_RDINS10(),
    .BRAM_RDINS11(),
    .BRAM_RDINS12(),
    .BRAM_RDINS13(),
    .BRAM_RDINS14(),
    .BRAM_RDINS15(),
    .BRAM_RDINS16(),
    .BRAM_RDINS17(),
    .BRAM_RDINS20(),
    .BRAM_RDINS24(),
    .BRAM_RDINS27(),
    .BRAM_RDINS28(),
    .BRAM_RDINS29(),
    .BRAM_RDINS31(),
    .BRAM_GCLKIN0(),
    .BRAM_GCLKIN1(\net_IBuf-clkpad-clk_BRAM_CLKH_VGCLK1_to_BRAM_GCLKIN15_1_0 ),
    .BRAM_GCLKIN2(),
    .BRAM_GCLKIN3(),
    .BRAM_GCLK_IOBD0(),
    .BRAM_GCLK_IOBD1(),
    .BRAM_GCLK_IOBD2(),
    .BRAM_GCLK_IOBD3(),
    .BRAM_GCLK_CLBD0(),
    .BRAM_GCLK_CLBD1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBD1_to_GCLK15_11_0 ),
    .BRAM_GCLK_CLBD2(),
    .BRAM_GCLK_CLBD3(),
    .BRAM_DIA6(),
    .BRAM_DIA7(),
    .BRAM_DIA14(),
    .BRAM_DIA15(),
    .BRAM_DIB6(),
    .BRAM_DIB7(),
    .BRAM_DIB14(),
    .BRAM_DIB15(),
    .BRAM_DOA3(),
    .BRAM_DOA7(),
    .BRAM_DOA11(),
    .BRAM_DOA15(),
    .BRAM_DOB3(),
    .BRAM_DOB7(),
    .BRAM_DOB11(),
    .BRAM_DOB15(),
    .BRAM_ADDRB8(),
    .BRAM_ADDRB9(),
    .BRAM_ADDRB10(),
    .BRAM_ADDRB11(),
    .BRAM_ADDRA8(),
    .BRAM_ADDRA9(),
    .BRAM_ADDRA10(),
    .BRAM_ADDRA11()
  );

  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufl0.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufl1.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufl2.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufl3.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufr0.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufr1.CONF = "0";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufr2.CONF = "1";
  defparam GSB_CLKV_5_28_0_inst.spbu_gclk_bufr3.CONF = "1";
  GSB_CLKV GSB_CLKV_5_28_0_inst (
    .CLKV_VGCLK0(),
    .CLKV_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK15_28_0 ),
    .CLKV_VGCLK2(),
    .CLKV_VGCLK3(),
    .CLKV_GCLK_BUFL0(),
    .CLKV_GCLK_BUFL1(),
    .CLKV_GCLK_BUFL2(),
    .CLKV_GCLK_BUFL3(),
    .CLKV_GCLK_BUFR0(),
    .CLKV_GCLK_BUFR1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFR1_to_GCLK15_32_0 ),
    .CLKV_GCLK_BUFR2(),
    .CLKV_GCLK_BUFR3()
  );

  defparam GSB_LBRAMC_4_1_0_inst.spbu_gclk_clbc0.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.spbu_gclk_clbc1.CONF = "0";
  defparam GSB_LBRAMC_4_1_0_inst.spbu_gclk_clbc2.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.spbu_gclk_clbc3.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.spbu_gclk_iobc0.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.spbu_gclk_iobc1.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.spbu_gclk_iobc2.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.spbu_gclk_iobc3.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.sps_addra4.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_addra5.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_addra6.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_addra7.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_addrb4.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_addrb5.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_addrb6.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_addrb7.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_clkb.CONF = "1111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_dia12.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_dia13.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_dia4.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_dia5.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_dib12.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_dib13.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_dib4.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_dib5.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec0.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec1.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec10.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec11.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec12.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec13.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec14.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec15.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec16.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec17.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec18.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec19.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec2.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec20.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec21.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec22.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec23.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec3.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec4.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec5.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec6.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec7.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec8.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_ec9.CONF = "11";
  defparam GSB_LBRAMC_4_1_0_inst.sps_h6bc0.CONF = "111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_h6bc1.CONF = "111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_h6bc2.CONF = "111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_h6bc3.CONF = "111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_h6mc0.CONF = "111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_h6mc1.CONF = "111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_h6mc2.CONF = "111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_h6mc3.CONF = "111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_lhc0.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_lhc3.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_lhc6.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_lhc9.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_llv1.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_llv5.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_llv9.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_raddrs1.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_raddrs13.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_raddrs17.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_raddrs21.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_raddrs25.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_raddrs29.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_raddrs5.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_raddrs9.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_rdins1.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_rdins13.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_rdins17.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_rdins21.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_rdins25.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_rdins29.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_rdins5.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_rdins9.CONF = "111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_rstb.CONF = "1111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_selb.CONF = "1111111";
  defparam GSB_LBRAMC_4_1_0_inst.sps_web.CONF = "1111111";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa10_rdouts10.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa10_rdouts27.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa14_rdouts12.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa14_rdouts29.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa2_rdouts10.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa2_rdouts27.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa2_rdouts28.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa2_rdouts9.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa6_rdouts11.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa6_rdouts12.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa6_rdouts29.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_doa6_rdouts30.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob10_rdouts11.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob10_rdouts28.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob14_rdouts13.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob14_rdouts30.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob2_rdouts10.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob2_rdouts11.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob2_rdouts28.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob2_rdouts29.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob6_rdouts12.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob6_rdouts13.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob6_rdouts30.CONF = "1";
  defparam GSB_LBRAMC_4_1_0_inst.tribuf_dob6_rdouts31.CONF = "1";
  GSB_LBRAMC GSB_LBRAMC_4_1_0_inst (
    .BRAM_EC0(),
    .BRAM_EC1(),
    .BRAM_EC2(),
    .BRAM_EC3(),
    .BRAM_EC4(),
    .BRAM_EC5(),
    .BRAM_EC6(),
    .BRAM_EC7(),
    .BRAM_EC8(),
    .BRAM_EC9(),
    .BRAM_EC10(),
    .BRAM_EC11(),
    .BRAM_EC12(),
    .BRAM_EC13(),
    .BRAM_EC14(),
    .BRAM_EC15(),
    .BRAM_EC16(),
    .BRAM_EC17(),
    .BRAM_EC18(),
    .BRAM_EC19(),
    .BRAM_EC20(),
    .BRAM_EC21(),
    .BRAM_EC22(),
    .BRAM_EC23(),
    .BRAM_H6EC0(),
    .BRAM_H6EC1(),
    .BRAM_H6EC2(),
    .BRAM_H6EC3(),
    .BRAM_H6BC0(),
    .BRAM_H6BC1(),
    .BRAM_H6BC2(),
    .BRAM_H6BC3(),
    .BRAM_H6MC0(),
    .BRAM_H6MC1(),
    .BRAM_H6MC2(),
    .BRAM_H6MC3(),
    .BRAM_H6DC0(),
    .BRAM_H6DC1(),
    .BRAM_H6DC2(),
    .BRAM_H6DC3(),
    .BRAM_LHC0(),
    .BRAM_LHC3(),
    .BRAM_LHC6(),
    .BRAM_LHC9(),
    .BRAM_LLV0(),
    .BRAM_LLV1(),
    .BRAM_LLV2(),
    .BRAM_LLV3(),
    .BRAM_LLV4(),
    .BRAM_LLV5(),
    .BRAM_LLV6(),
    .BRAM_LLV7(),
    .BRAM_LLV8(),
    .BRAM_LLV9(),
    .BRAM_LLV10(),
    .BRAM_LLV11(),
    .BRAM_RDOUTS1(),
    .BRAM_RDOUTS5(),
    .BRAM_RDOUTS9(),
    .BRAM_RDOUTS10(),
    .BRAM_RDOUTS11(),
    .BRAM_RDOUTS12(),
    .BRAM_RDOUTS13(),
    .BRAM_RDOUTS17(),
    .BRAM_RDOUTS21(),
    .BRAM_RDOUTS25(),
    .BRAM_RDOUTS27(),
    .BRAM_RDOUTS28(),
    .BRAM_RDOUTS29(),
    .BRAM_RDOUTS30(),
    .BRAM_RDOUTS31(),
    .BRAM_RDINS1(),
    .BRAM_RDINS2(),
    .BRAM_RDINS3(),
    .BRAM_RDINS5(),
    .BRAM_RDINS6(),
    .BRAM_RDINS7(),
    .BRAM_RDINS9(),
    .BRAM_RDINS13(),
    .BRAM_RDINS17(),
    .BRAM_RDINS19(),
    .BRAM_RDINS20(),
    .BRAM_RDINS21(),
    .BRAM_RDINS23(),
    .BRAM_RDINS24(),
    .BRAM_RDINS25(),
    .BRAM_RDINS29(),
    .BRAM_RADDRS0(),
    .BRAM_RADDRS1(),
    .BRAM_RADDRS2(),
    .BRAM_RADDRS3(),
    .BRAM_RADDRS5(),
    .BRAM_RADDRS8(),
    .BRAM_RADDRS9(),
    .BRAM_RADDRS10(),
    .BRAM_RADDRS11(),
    .BRAM_RADDRS12(),
    .BRAM_RADDRS13(),
    .BRAM_RADDRS14(),
    .BRAM_RADDRS15(),
    .BRAM_RADDRS16(),
    .BRAM_RADDRS17(),
    .BRAM_RADDRS18(),
    .BRAM_RADDRS19(),
    .BRAM_RADDRS21(),
    .BRAM_RADDRS24(),
    .BRAM_RADDRS25(),
    .BRAM_RADDRS26(),
    .BRAM_RADDRS27(),
    .BRAM_RADDRS28(),
    .BRAM_RADDRS29(),
    .BRAM_RADDRS30(),
    .BRAM_RADDRS31(),
    .BRAM_DIA4(),
    .BRAM_DIA5(),
    .BRAM_DIA12(),
    .BRAM_DIA13(),
    .BRAM_DIB4(),
    .BRAM_DIB5(),
    .BRAM_DIB12(),
    .BRAM_DIB13(),
    .BRAM_DOA2(),
    .BRAM_DOA6(),
    .BRAM_DOA10(),
    .BRAM_DOA14(),
    .BRAM_DOB2(),
    .BRAM_DOB6(),
    .BRAM_DOB10(),
    .BRAM_DOB14(),
    .BRAM_ADDRA4(),
    .BRAM_ADDRA5(),
    .BRAM_ADDRA6(),
    .BRAM_ADDRA7(),
    .BRAM_ADDRB4(),
    .BRAM_ADDRB5(),
    .BRAM_ADDRB6(),
    .BRAM_ADDRB7(),
    .BRAM_CLKB(),
    .BRAM_WEB(),
    .BRAM_SELB(),
    .BRAM_RSTB(),
    .BRAM_GCLKIN0(),
    .BRAM_GCLKIN1(\net_IBuf-clkpad-clk_BRAM_CLKH_VGCLK1_to_BRAM_GCLKIN15_1_0 ),
    .BRAM_GCLKIN2(),
    .BRAM_GCLKIN3(),
    .BRAM_GCLK_IOBC0(),
    .BRAM_GCLK_IOBC1(),
    .BRAM_GCLK_IOBC2(),
    .BRAM_GCLK_IOBC3(),
    .BRAM_GCLK_CLBC0(),
    .BRAM_GCLK_CLBC1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBC1_to_GCLK14_11_0 ),
    .BRAM_GCLK_CLBC2(),
    .BRAM_GCLK_CLBC3()
  );

  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufl0.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufl1.CONF = "0";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufl2.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufl3.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufr0.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufr1.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufr2.CONF = "1";
  defparam GSB_CLKV_6_28_0_inst.spbu_gclk_bufr3.CONF = "1";
  GSB_CLKV GSB_CLKV_6_28_0_inst (
    .CLKV_VGCLK0(),
    .CLKV_VGCLK1(\net_IBuf-clkpad-clk_CLKC_VGCLK1_to_CLKV_VGCLK15_28_0 ),
    .CLKV_VGCLK2(),
    .CLKV_VGCLK3(),
    .CLKV_GCLK_BUFL0(),
    .CLKV_GCLK_BUFL1(\net_IBuf-clkpad-clk_CLKV_GCLK_BUFL1_to_GCLK16_16_0 ),
    .CLKV_GCLK_BUFL2(),
    .CLKV_GCLK_BUFL3(),
    .CLKV_GCLK_BUFR0(),
    .CLKV_GCLK_BUFR1(),
    .CLKV_GCLK_BUFR2(),
    .CLKV_GCLK_BUFR3()
  );

  defparam GSB_CNT_3_40_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_h6w2.CONF = "0010";
  defparam GSB_CNT_3_40_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_40_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_40_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_out7.CONF = "101101";
  defparam GSB_CNT_3_40_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e1.CONF = "01";
  defparam GSB_CNT_3_40_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e11.CONF = "01";
  defparam GSB_CNT_3_40_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_e20.CONF = "0";
  defparam GSB_CNT_3_40_0_inst.sps_e21.CONF = "01";
  defparam GSB_CNT_3_40_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_out1.CONF = "000111";
  defparam GSB_CNT_3_40_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_out3.CONF = "000111";
  defparam GSB_CNT_3_40_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_out5.CONF = "011110";
  defparam GSB_CNT_3_40_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_s0_bx_b.CONF = "011011";
  defparam GSB_CNT_3_40_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_f_b1.CONF = "001101111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_f_b2.CONF = "010101111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_s1_bx_b.CONF = "001101";
  defparam GSB_CNT_3_40_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s1_f_b1.CONF = "010101111";
  defparam GSB_CNT_3_40_0_inst.sps_s1_f_b2.CONF = "001111101";
  defparam GSB_CNT_3_40_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_40_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_40_0_inst.sps_s1_g_b1.CONF = "010011";
  defparam GSB_CNT_3_40_0_inst.sps_s1_g_b2.CONF = "001100";
  defparam GSB_CNT_3_40_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_s2.CONF = "01";
  defparam GSB_CNT_3_40_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_40_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_40_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_40_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_40_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e17_w17.CONF = "0";
  defparam GSB_CNT_3_40_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e3_w3.CONF = "0";
  defparam GSB_CNT_3_40_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_40_0_inst.switch_s9_n9.CONF = "0";
  defparam GSB_CNT_3_40_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_40_0_inst (
    .E0(),
    .E1(\net_Buf-pad-RGB[12]_E1_to_W13_42_0 ),
    .E2(),
    .E3(\net_Buf-pad-RGB[23]_W3_to_E33_40_0 ),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(net_U9_CO_W10_to_E103_40_0),
    .E11(net_U14_S_E11_to_W113_42_0),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(net_U10_S_E17_to_W173_42_0),
    .E18(),
    .E19(),
    .E20(net_U8_CO_E20_to_W203_42_0),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(\net_Buf-pad-RGB[22]_S9_to_N93_40_0 ),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(\net_Buf-pad-RGB[6]_S16_to_N163_40_0 ),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(\net_Buf-pad-RGB[22]_S21_to_N213_40_0 ),
    .N22(\net_Buf-pad-RGB[13]_S22_to_N223_40_0 ),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(\net_Buf-pad-RGB[23]_W3_to_E33_39_0 ),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(net_U10_S_E14_to_W143_40_0),
    .W15(),
    .W16(),
    .W17(net_U10_S_E17_to_W173_40_0),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(net_U7_S_H6W2_to_H6E23_34_0),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(net_U14_S_OUT1_to_OUT_W13_42_0),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(\net_Buf-pad-RGB[13]_TOP_V6B0_to_V6N03_40_0 ),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(\net_Buf-pad-RGB[12]_TOP_V6D0_to_V6M03_40_0 ),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(\net_Buf-pad-RGB[6]_TOP_V6D10_to_V6M103_40_0 ),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-RGB[13]_S0_F_B1_to_F13_40_0 ),
    .S0_F_B2(\net_Buf-pad-RGB[6]_S0_F_B2_to_F23_40_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(\net_Buf-pad-RGB[22]_S0_BX_B_to_BX3_40_0 ),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(net_U14_S_X_to_S0_X3_40_0),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Buf-pad-RGB[13]_S1_F_B1_to_F13_40_0 ),
    .S1_F_B2(\net_Buf-pad-RGB[6]_S1_F_B2_to_F23_40_0 ),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(net_U10_S_S1_G_B1_to_G13_40_0),
    .S1_G_B2(net_U9_CO_S1_G_B2_to_G23_40_0),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(\net_Buf-pad-RGB[22]_S1_BX_B_to_BX3_40_0 ),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(net_U8_CO_XB_to_S1_XB3_40_0),
    .S1_Y(net_U7_S_Y_to_S1_Y3_40_0),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_3_34_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_h6w2.CONF = "0000";
  defparam GSB_CNT_3_34_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_34_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_34_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_e21.CONF = "01";
  defparam GSB_CNT_3_34_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_e9.CONF = "01";
  defparam GSB_CNT_3_34_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_34_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_34_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_34_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_34_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_34_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_34_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(\net_Buf-pad-RGB[15]_E9_to_W93_35_0 ),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(\net_Buf-pad-RGB[15]_E21_to_W213_35_0 ),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(net_U7_S_H6W2_to_H6E23_34_0),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(net_U7_S_H6W2_to_H6M23_31_0),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(\net_Buf-pad-RGB[15]_TOP_V6D8_to_V6M83_34_0 ),
    .V6M9(),
    .V6M10(\net_Buf-pad-RGB[15]_TOP_V6D10_to_V6M103_34_0 ),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_3_31_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_31_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_31_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_v6s2.CONF = "0011";
  defparam GSB_CNT_3_31_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_31_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_31_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_31_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_31_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_31_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_31_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(net_U7_S_H6W2_to_H6M23_31_0),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(net_U7_S_V6S2_to_V6M26_31_0),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_31_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_31_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_31_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e13.CONF = "01";
  defparam GSB_CNT_6_31_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_31_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_31_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_31_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_31_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_31_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_31_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(net_U7_S_E13_to_W136_32_0),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(net_U7_S_V6S2_to_V6M26_31_0),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_32_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_32_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_32_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_32_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_32_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_32_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_32_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n8_w13.CONF = "0";
  defparam GSB_CNT_6_32_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_32_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_32_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(net_U7_S_N8_to_S85_32_0),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(net_U7_S_E13_to_W136_32_0),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_3_42_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_h6w10.CONF = "000";
  defparam GSB_CNT_3_42_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_h6w4.CONF = "000";
  defparam GSB_CNT_3_42_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_h6w8.CONF = "101";
  defparam GSB_CNT_3_42_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_42_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_42_0_inst.sps_out6.CONF = "011011";
  defparam GSB_CNT_3_42_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_w10.CONF = "10";
  defparam GSB_CNT_3_42_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w3.CONF = "10";
  defparam GSB_CNT_3_42_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_n12.CONF = "01";
  defparam GSB_CNT_3_42_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_out0.CONF = "011110";
  defparam GSB_CNT_3_42_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_out3.CONF = "010111";
  defparam GSB_CNT_3_42_0_inst.sps_out4.CONF = "101101";
  defparam GSB_CNT_3_42_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s0_f_b1.CONF = "110111111";
  defparam GSB_CNT_3_42_0_inst.sps_s0_f_b2.CONF = "010110111";
  defparam GSB_CNT_3_42_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_42_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_42_0_inst.sps_s0_g_b1.CONF = "100010";
  defparam GSB_CNT_3_42_0_inst.sps_s0_g_b2.CONF = "010011";
  defparam GSB_CNT_3_42_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s15.CONF = "01";
  defparam GSB_CNT_3_42_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_s1_bx_b.CONF = "000111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_f_b1.CONF = "100101111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_f_b2.CONF = "100110111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_g_b1.CONF = "001111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_g_b2.CONF = "100000";
  defparam GSB_CNT_3_42_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_42_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_42_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_42_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_42_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s9_e11.CONF = "0";
  defparam GSB_CNT_3_42_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_42_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_42_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(net_U18_S_W11_to_E113_42_0),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(\net_Buf-pad-RGB[5]_S2_to_N23_42_0 ),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(\net_Buf-pad-RGB[21]_S15_to_N153_42_0 ),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(\net_Buf-pad-RGB[12]_E1_to_W13_42_0 ),
    .W2(),
    .W3(\net_Buf-pad-RGB[23]_W3_to_E33_40_0 ),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(net_U9_CO_W10_to_E103_40_0),
    .W11(net_U14_S_E11_to_W113_42_0),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(net_U10_S_E17_to_W173_42_0),
    .W18(),
    .W19(),
    .W20(net_U8_CO_E20_to_W203_42_0),
    .W21(),
    .W22(),
    .W23(),
    .S0(net_U13_CO_boy_net_N0_to_S03_42_0),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(net_U18_S_S9_to_N94_42_0),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(\net_Buf-pad-RGB[20]_S15_to_N154_42_0 ),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(\net_Buf-pad-RGB[23]_H6W4_to_H6E43_42_0 ),
    .H6E5(),
    .H6E6(\net_Buf-pad-RGB[20]_H6W6_to_H6E63_42_0 ),
    .H6E7(),
    .H6E8(\net_Buf-pad-RGB[23]_H6W8_to_H6E83_42_0 ),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(net_U11_S_H6W4_to_H6E43_35_0),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(\net_Buf-pad-RGB[23]_H6W8_to_H6E83_35_0 ),
    .H6W9(),
    .H6W10(net_U6_CO_H6W10_to_H6E103_35_0),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(net_U14_S_OUT1_to_OUT_W13_42_0),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(net_U14_S_S0_F_B1_to_F13_42_0),
    .S0_F_B2(net_U12_CO_S0_F_B2_to_F23_42_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(net_U10_S_S0_G_B1_to_G13_42_0),
    .S0_G_B2(net_U8_CO_S0_G_B2_to_G23_42_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(net_U9_CO_XB_to_S0_XB3_42_0),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(net_U6_CO_COUT_to_CO_0_LOCAL3_42_0),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Buf-pad-RGB[12]_S1_F_B1_to_F13_42_0 ),
    .S1_F_B2(\net_Buf-pad-RGB[5]_S1_F_B2_to_F23_42_0 ),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(net_U14_S_S1_G_B1_to_G13_42_0),
    .S1_G_B2(net_U13_CO_boy_net_S1_G_B2_to_G23_42_0),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(\net_Buf-pad-RGB[21]_S1_BX_B_to_BX3_42_0 ),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(net_U12_CO_XB_to_S1_XB3_42_0),
    .S1_Y(net_U11_S_Y_to_S1_Y3_42_0),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_3_32_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_32_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_32_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_s2.CONF = "10";
  defparam GSB_CNT_3_32_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_32_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_32_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_32_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_32_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_32_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_32_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(net_U11_S_S2_to_N24_32_0),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(net_U11_S_H6W4_to_H6M43_32_0),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_32_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_32_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_32_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_32_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_32_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_32_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_32_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s2_n2.CONF = "0";
  defparam GSB_CNT_4_32_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_32_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_32_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(net_U11_S_S2_to_N24_32_0),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(net_U11_S_S2_to_N25_32_0),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_42_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_llh0.CONF = "01";
  defparam GSB_CNT_4_42_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_42_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_42_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_e7.CONF = "0";
  defparam GSB_CNT_4_42_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_h6e2.CONF = "0011";
  defparam GSB_CNT_4_42_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_n0.CONF = "01";
  defparam GSB_CNT_4_42_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n13.CONF = "10";
  defparam GSB_CNT_4_42_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_out0.CONF = "011011";
  defparam GSB_CNT_4_42_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_out2.CONF = "101101";
  defparam GSB_CNT_4_42_0_inst.sps_out3.CONF = "011110";
  defparam GSB_CNT_4_42_0_inst.sps_out4.CONF = "010111";
  defparam GSB_CNT_4_42_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_s0_bx_b.CONF = "001011";
  defparam GSB_CNT_4_42_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s0_f_b1.CONF = "100111011";
  defparam GSB_CNT_4_42_0_inst.sps_s0_f_b2.CONF = "001111101";
  defparam GSB_CNT_4_42_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_42_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_42_0_inst.sps_s0_g_b1.CONF = "011000";
  defparam GSB_CNT_4_42_0_inst.sps_s0_g_b2.CONF = "001101";
  defparam GSB_CNT_4_42_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s16.CONF = "01";
  defparam GSB_CNT_4_42_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_s1_bx_b.CONF = "000111";
  defparam GSB_CNT_4_42_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s1_f_b1.CONF = "100111101";
  defparam GSB_CNT_4_42_0_inst.sps_s1_f_b2.CONF = "011110111";
  defparam GSB_CNT_4_42_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_42_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_42_0_inst.sps_s1_g_b1.CONF = "011111";
  defparam GSB_CNT_4_42_0_inst.sps_s1_g_b2.CONF = "011011";
  defparam GSB_CNT_4_42_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s7.CONF = "0";
  defparam GSB_CNT_4_42_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_42_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_42_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_42_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_42_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n11_w12.CONF = "0";
  defparam GSB_CNT_4_42_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n14_e10.CONF = "0";
  defparam GSB_CNT_4_42_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_42_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_42_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(\net_Buf-pad-RGB[11]_E7_to_W74_43_0 ),
    .E8(net_U18_S_W8_to_E84_42_0),
    .E9(),
    .E10(net_U23_S_W10_to_E104_42_0),
    .E11(\net_Lut-U21_0_0_W11_to_E114_42_0 ),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(net_U13_CO_boy_net_N0_to_S03_42_0),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(net_U18_S_S9_to_N94_42_0),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(\net_Buf-pad-RGB[20]_S15_to_N154_42_0 ),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(net_U20_CO_E4_to_W44_42_0),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_Buf-pad-RGB[4]_E12_to_W124_42_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(net_U15_S_LLH0_to_LLH64_9_0),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(\net_Buf-pad-RGB[11]_TOP_V6M2_to_V6N24_42_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_Buf-pad-RGB[11]_TOP_V6S1_to_V6M14_42_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(net_U23_S_S0_F_B1_to_F14_42_0),
    .S0_F_B2(\net_Lut-U21_0_0_S0_F_B2_to_F24_42_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(net_U18_S_S0_G_B1_to_G14_42_0),
    .S0_G_B2(net_U16_CO_S0_G_B2_to_G24_42_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(net_U20_CO_S0_BX_B_to_BX4_42_0),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(net_U17_CO_XB_to_S0_XB4_42_0),
    .S0_Y(),
    .S0_YB(net_U13_CO_boy_net_YB_to_S0_YB4_42_0),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(net_U13_CO_COUT_to_CO_0_LOCAL4_42_0),
    .CO_0(net_U13_CO_CO_0_to_CIN4_42_0),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Buf-pad-RGB[11]_S1_F_B1_to_F14_42_0 ),
    .S1_F_B2(\net_Buf-pad-RGB[4]_S1_F_B2_to_F24_42_0 ),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(net_U18_S_S1_G_B1_to_G14_42_0),
    .S1_G_B2(net_U17_CO_S1_G_B2_to_G24_42_0),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(\net_Buf-pad-RGB[20]_S1_BX_B_to_BX4_42_0 ),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(net_U16_CO_XB_to_S1_XB4_42_0),
    .S1_Y(net_U15_S_Y_to_S1_Y4_42_0),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_9_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_9_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_9_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_h6e3.CONF = "0001";
  defparam GSB_CNT_4_9_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_9_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_9_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_9_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_9_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_9_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_9_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(net_U15_S_H6E3_to_H6M34_12_0),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(net_U15_S_LLH0_to_LLH64_9_0),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_12_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_12_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_12_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s21.CONF = "0";
  defparam GSB_CNT_4_12_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_12_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_12_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_12_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_12_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s21_w3.CONF = "0";
  defparam GSB_CNT_4_12_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_12_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_12_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(net_U15_S_W3_to_E34_11_0),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(net_U15_S_H6E3_to_H6M34_12_0),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_44_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_4_44_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_44_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_44_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w11.CONF = "01";
  defparam GSB_CNT_4_44_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_w15.CONF = "10";
  defparam GSB_CNT_4_44_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_n18.CONF = "01";
  defparam GSB_CNT_4_44_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_out5.CONF = "000111";
  defparam GSB_CNT_4_44_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_f_b1.CONF = "110111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_f_b2.CONF = "100110111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s10.CONF = "01";
  defparam GSB_CNT_4_44_0_inst.sps_s11.CONF = "0";
  defparam GSB_CNT_4_44_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s14.CONF = "01";
  defparam GSB_CNT_4_44_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_44_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_44_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_44_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_44_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_44_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_44_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(\net_Lut-U21_0_0_W11_to_E114_43_0 ),
    .W12(),
    .W13(),
    .W14(),
    .W15(\net_Buf-pad-RGB[4]_W15_to_E154_43_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(\net_Buf-pad-RGB[10]_S10_to_N105_44_0 ),
    .S11(\net_Buf-pad-RGB[9]_S11_to_N115_44_0 ),
    .S12(),
    .S13(),
    .S14(\net_Buf-pad-RGB[10]_S14_to_N145_44_0 ),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(\net_Lut-U21_0_0_H6W3_to_H6E34_44_0 ),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(\net_Lut-U21_0_0_H6W8_to_H6E84_44_0 ),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(\net_Buf-pad-RGB[9]_H6W8_to_H6M84_44_0 ),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(net_U19_S_LLH6_to_LLH04_11_0),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(net_U23_S_OUT1_to_OUT_W14_44_0),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(\net_Buf-pad-RGB[10]_TOP_V6M1_to_V6N14_44_0 ),
    .V6N2(\net_Buf-pad-RGB[10]_TOP_V6M2_to_V6N24_44_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(\net_Buf-pad-RGB[4]_TOP_V6S2_to_V6M24_44_0 ),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(net_U23_S_S0_F_B1_to_F14_44_0),
    .S0_F_B2(\net_Lut-U21_0_0_S0_F_B2_to_F24_44_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(net_U19_S_X_to_S0_X4_44_0),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_44_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_h6w1.CONF = "0010";
  defparam GSB_CNT_5_44_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_llh6.CONF = "01";
  defparam GSB_CNT_5_44_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_44_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_44_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_e6.CONF = "10";
  defparam GSB_CNT_5_44_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_out2.CONF = "010111";
  defparam GSB_CNT_5_44_0_inst.sps_out3.CONF = "011011";
  defparam GSB_CNT_5_44_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_out5.CONF = "011101";
  defparam GSB_CNT_5_44_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_s0_bx_b.CONF = "001101";
  defparam GSB_CNT_5_44_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s0_f_b1.CONF = "011111101";
  defparam GSB_CNT_5_44_0_inst.sps_s0_f_b2.CONF = "001101111";
  defparam GSB_CNT_5_44_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_44_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_44_0_inst.sps_s0_g_b1.CONF = "100101";
  defparam GSB_CNT_5_44_0_inst.sps_s0_g_b2.CONF = "010101";
  defparam GSB_CNT_5_44_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s14.CONF = "10";
  defparam GSB_CNT_5_44_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_s1_bx_b.CONF = "111110";
  defparam GSB_CNT_5_44_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s1_f_b1.CONF = "010111011";
  defparam GSB_CNT_5_44_0_inst.sps_s1_f_b2.CONF = "010111011";
  defparam GSB_CNT_5_44_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_44_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_44_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s23.CONF = "0";
  defparam GSB_CNT_5_44_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_44_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_44_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_44_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_44_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_44_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_44_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(\net_Buf-pad-RGB[10]_S10_to_N105_44_0 ),
    .N11(\net_Buf-pad-RGB[9]_S11_to_N115_44_0 ),
    .N12(),
    .N13(),
    .N14(\net_Buf-pad-RGB[10]_S14_to_N145_44_0 ),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(\net_Buf-pad-RGB[18]_E13_to_W135_44_0 ),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(\net_Buf-pad-RGB[2]_N19_to_S195_44_0 ),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(\net_Lut-U26_0InvLut_H6W6_to_H6M65_44_0 ),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(\net_Lut-U26_0InvLut_H6W10_to_H6M105_44_0 ),
    .H6M11(),
    .H6W0(),
    .H6W1(net_U20_CO_H6W1_to_H6M15_40_0),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(net_U24_S_LLH6_to_LLH65_18_0),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-RGB[18]_S0_F_B1_to_F15_44_0 ),
    .S0_F_B2(\net_Buf-pad-RGB[2]_S0_F_B2_to_F25_44_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Buf-pad-RGB[10]_S0_G_B1_to_G15_44_0 ),
    .S0_G_B2(\net_Lut-U26_0InvLut_S0_G_B2_to_G25_44_0 ),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(\net_Buf-pad-RGB[9]_S0_BX_B_to_BX5_44_0 ),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(net_U25_CO_XB_to_S0_XB5_44_0),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(net_U20_CO_COUT_to_CO_0_LOCAL5_44_0),
    .CO_0(net_U20_CO_CO_0_to_CIN5_44_0),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Buf-pad-RGB[10]_S1_F_B1_to_F15_44_0 ),
    .S1_F_B2(\net_Lut-U26_0InvLut_S1_F_B2_to_F25_44_0 ),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(net_U25_CO_S1_BX_B_to_BX5_44_0),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(net_U24_S_X_to_S1_X5_44_0),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_18_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w2.CONF = "0001";
  defparam GSB_CNT_5_18_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_18_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_18_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_18_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_18_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_18_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_18_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_18_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(net_U24_S_H6W2_to_H6M25_14_0),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(net_U24_S_LLH6_to_LLH65_18_0),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_14_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_14_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_14_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s18.CONF = "10";
  defparam GSB_CNT_5_14_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_14_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_14_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_14_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_14_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_14_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(net_U24_S_S18_to_N186_14_0),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(net_U24_S_H6W2_to_H6M25_14_0),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_14_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_14_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_14_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_14_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_14_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_14_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_14_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n18_e14.CONF = "0";
  defparam GSB_CNT_6_14_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_14_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_14_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(net_U24_S_E14_to_W146_16_0),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(net_U24_S_S18_to_N186_14_0),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_45_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_llh0.CONF = "01";
  defparam GSB_CNT_5_45_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_45_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_45_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_out3.CONF = "000111";
  defparam GSB_CNT_5_45_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_s0_bx_b.CONF = "111101";
  defparam GSB_CNT_5_45_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s0_f_b1.CONF = "011111011";
  defparam GSB_CNT_5_45_0_inst.sps_s0_f_b2.CONF = "001111110";
  defparam GSB_CNT_5_45_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_45_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_45_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s6.CONF = "10";
  defparam GSB_CNT_5_45_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_45_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_45_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_45_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_45_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_45_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_45_0_inst (
    .E0(),
    .E1(\net_Buf-pad-RGB[9]_W1_to_E15_45_0 ),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(\net_Buf-pad-RGB[2]_N4_to_S45_45_0 ),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(\net_Buf-pad-RGB[18]_H6W0_to_H6M05_45_0 ),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(net_U27_S_LLH0_to_LLH05_19_0),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-RGB[18]_S0_F_B1_to_F15_45_0 ),
    .S0_F_B2(\net_Buf-pad-RGB[2]_S0_F_B2_to_F25_45_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(\net_Buf-pad-RGB[9]_S0_BX_B_to_BX5_45_0 ),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(net_U27_S_X_to_S0_X5_45_0),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_16_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_16_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_16_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s6.CONF = "10";
  defparam GSB_CNT_5_16_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_16_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_16_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_16_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_16_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_16_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_16_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(net_U27_S_S6_to_N66_16_0),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(net_U27_S_H6W0_to_H6M05_16_0),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_21_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_21_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_21_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6e1.CONF = "01011011";
  defparam GSB_TOP_1_21_0_inst.sps_h6e2.CONF = "01011011";
  defparam GSB_TOP_1_21_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_21_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_21_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_21_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_21_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_21_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(\net_Buf-pad-RGB[15]_TOP_H6E1_to_TOP_H6W11_27_0 ),
    .TOP_H6E2(\net_Buf-pad-RGB[15]_TOP_H6E2_to_TOP_H6W21_27_0 ),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(\net_Buf-pad-RGB[15]_IN_to_TOP_I11_21_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_27_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_27_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_27_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6e1.CONF = "01101110";
  defparam GSB_TOP_1_27_0_inst.sps_h6e2.CONF = "01101110";
  defparam GSB_TOP_1_27_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_27_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_27_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_27_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_27_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_27_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(\net_Buf-pad-RGB[15]_TOP_H6E1_to_TOP_H6W11_34_0 ),
    .TOP_H6E2(\net_Buf-pad-RGB[15]_TOP_H6E2_to_TOP_H6W21_34_0 ),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(\net_Buf-pad-RGB[15]_TOP_H6E1_to_TOP_H6W11_27_0 ),
    .TOP_H6W2(\net_Buf-pad-RGB[15]_TOP_H6E2_to_TOP_H6W21_27_0 ),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_34_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_34_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_34_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_34_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_34_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d10.CONF = "111011";
  defparam GSB_TOP_1_34_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_34_0_inst.sps_v6d8.CONF = "111011";
  defparam GSB_TOP_1_34_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_34_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_34_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(\net_Buf-pad-RGB[15]_TOP_H6E1_to_TOP_H6W11_34_0 ),
    .TOP_H6W2(\net_Buf-pad-RGB[15]_TOP_H6E2_to_TOP_H6W21_34_0 ),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(\net_Buf-pad-RGB[15]_TOP_V6D8_to_V6M83_34_0 ),
    .TOP_V6D9(),
    .TOP_V6D10(\net_Buf-pad-RGB[15]_TOP_V6D10_to_V6M103_34_0 ),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_35_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_35_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_35_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6e2.CONF = "01011011";
  defparam GSB_TOP_1_35_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_35_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_35_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d0.CONF = "01101";
  defparam GSB_TOP_1_35_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d10.CONF = "101111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_35_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_35_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_35_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(\net_Buf-pad-RGB[14]_TOP_H6E2_to_TOP_H6M21_38_0 ),
    .TOP_H6E3(\net_Buf-pad-RGB[7]_TOP_H6W3_to_TOP_H6E31_35_0 ),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(\net_Buf-pad-RGB[14]_TOP_V6D0_to_V6M03_35_0 ),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(\net_Buf-pad-RGB[7]_TOP_V6D10_to_V6M103_35_0 ),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(\net_Buf-pad-RGB[14]_IN_to_TOP_I11_35_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_38_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_38_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_38_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_38_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_38_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_38_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_38_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_38_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6d10.CONF = "110111";
  defparam GSB_TOP_1_38_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_v6d6.CONF = "110111";
  defparam GSB_TOP_1_38_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_38_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_38_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_38_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(\net_Buf-pad-RGB[7]_TOP_H6W0_to_TOP_H6M01_38_0 ),
    .TOP_H6M1(),
    .TOP_H6M2(\net_Buf-pad-RGB[14]_TOP_H6E2_to_TOP_H6M21_38_0 ),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(\net_Buf-pad-RGB[7]_TOP_V6D6_to_V6M63_38_0 ),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(\net_Buf-pad-RGB[14]_TOP_V6D10_to_V6M103_38_0 ),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_CNT_3_38_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_38_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_38_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e12.CONF = "10";
  defparam GSB_CNT_3_38_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_e21.CONF = "01";
  defparam GSB_CNT_3_38_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_38_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_38_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_38_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_38_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_38_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_38_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(\net_Buf-pad-RGB[7]_E12_to_W123_39_0 ),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(\net_Buf-pad-RGB[14]_E21_to_W213_39_0 ),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(\net_Buf-pad-RGB[7]_TOP_V6D6_to_V6M63_38_0 ),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(\net_Buf-pad-RGB[14]_TOP_V6D10_to_V6M103_38_0 ),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_3_39_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_39_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_39_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e14.CONF = "0";
  defparam GSB_CNT_3_39_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_e17.CONF = "10";
  defparam GSB_CNT_3_39_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_out4.CONF = "000111";
  defparam GSB_CNT_3_39_0_inst.sps_out5.CONF = "000111";
  defparam GSB_CNT_3_39_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_s0_bx_b.CONF = "011101";
  defparam GSB_CNT_3_39_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_f_b1.CONF = "010101111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_f_b2.CONF = "001110111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_39_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_39_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_39_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_39_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_39_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_39_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(\net_Buf-pad-RGB[23]_W3_to_E33_39_0 ),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(net_U10_S_E14_to_W143_40_0),
    .E15(),
    .E16(),
    .E17(net_U10_S_E17_to_W173_40_0),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_Buf-pad-RGB[7]_E12_to_W123_39_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(\net_Buf-pad-RGB[14]_E21_to_W213_39_0 ),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-RGB[14]_S0_F_B1_to_F13_39_0 ),
    .S0_F_B2(\net_Buf-pad-RGB[7]_S0_F_B2_to_F23_39_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(\net_Buf-pad-RGB[23]_S0_BX_B_to_BX3_39_0 ),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(net_U10_S_X_to_S0_X3_39_0),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_48_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6w0.CONF = "01011110";
  defparam GSB_TOP_1_48_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6w3.CONF = "01011110";
  defparam GSB_TOP_1_48_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_48_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_48_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_48_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_48_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_48_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_48_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_48_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(\net_Buf-pad-RGB[7]_TOP_H6W0_to_TOP_H6E01_42_0 ),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(\net_Buf-pad-RGB[7]_TOP_H6W3_to_TOP_H6E31_42_0 ),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(\net_Buf-pad-RGB[7]_IN_to_TOP_I21_48_0 ),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_42_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6w0.CONF = "01101110";
  defparam GSB_TOP_1_42_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6w3.CONF = "01101110";
  defparam GSB_TOP_1_42_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_42_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_42_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s1.CONF = "0111110";
  defparam GSB_TOP_1_42_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_42_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv11.CONF = "00";
  defparam GSB_TOP_1_42_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_42_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_42_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_42_0_inst.sps_v6m2.CONF = "01101";
  defparam GSB_TOP_1_42_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_42_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(\net_Buf-pad-RGB[7]_TOP_H6W0_to_TOP_H6E01_42_0 ),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(\net_Buf-pad-RGB[7]_TOP_H6W3_to_TOP_H6E31_42_0 ),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(\net_Buf-pad-RGB[5]_TOP_H6W4_to_TOP_H6A41_42_0 ),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(\net_Buf-pad-RGB[7]_TOP_H6W0_to_TOP_H6M01_38_0 ),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(\net_Buf-pad-RGB[7]_TOP_H6W3_to_TOP_H6E31_35_0 ),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(\net_Buf-pad-RGB[11]_TOP_V6M2_to_V6N24_42_0 ),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(\net_Buf-pad-RGB[11]_TOP_V6S1_to_V6M14_42_0 ),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(\net_Buf-pad-RGB[5]_TOP_LLV11_to_LLV02_42_0 ),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(\net_Buf-pad-RGB[11]_IN_to_TOP_I21_42_0 ),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_RHT_34_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_34_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_34_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_34_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_34_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_34_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_34_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_34_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_34_54_0_inst.sps_llv6.CONF = "0011011111";
  defparam GSB_RHT_34_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_34_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_34_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_34_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_34_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_34_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_34_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_34_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_34_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_34_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_34_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_34_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_34_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_34_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_34_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_34_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_34_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(),
    .RIGHT_LLV6(\net_Buf-pad-RGB[23]_RIGHT_LLV6_to_RIGHT_LLV03_54_0 ),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(\net_Buf-pad-RGB[23]_IN_to_RIGHT_I234_54_0 ),
    .RIGHT_I3(),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_RHT_3_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_3_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_3_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_3_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_3_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_3_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_3_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_3_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_3_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6d4.CONF = "101111";
  defparam GSB_RHT_3_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_3_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_3_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_3_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_3_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_h6w4.CONF = "111011";
  defparam GSB_RHT_3_54_0_inst.sps_h6w6.CONF = "111011";
  defparam GSB_RHT_3_54_0_inst.sps_h6w8.CONF = "101111";
  defparam GSB_RHT_3_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_3_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_3_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_3_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_3_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_3_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_3_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_3_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_3_54_0_inst.sps_v6n0.CONF = "00111011";
  defparam GSB_RHT_3_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_3_54_0_inst.sps_v6n2.CONF = "00111011";
  defparam GSB_RHT_3_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_3_54_0_inst.sps_v6s0.CONF = "00111011";
  defparam GSB_RHT_3_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_3_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_3_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_3_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_3_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_3_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_3_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_3_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_3_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_3_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_3_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_3_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_3_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(\net_Buf-pad-RGB[20]_RIGHT_H6D4_to_H6E43_49_0 ),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(\net_Buf-pad-RGB[23]_RIGHT_H6W4_to_H6E43_48_0 ),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(\net_Buf-pad-RGB[20]_RIGHT_H6W6_to_H6E63_48_0 ),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(\net_Buf-pad-RGB[23]_RIGHT_H6W8_to_H6E83_48_0 ),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(\net_Buf-pad-RGB[20]_UR_V6B1_to_RIGHT_V6N13_54_0 ),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(\net_Buf-pad-RGB[23]_RIGHT_LLV6_to_RIGHT_LLV03_54_0 ),
    .RIGHT_LLV6(\net_Buf-pad-RGB[20]_RIGHT_LLV6_to_UR_LLV41_54_0 ),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(),
    .RIGHT_I3(),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_3_48_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_h6w4.CONF = "101";
  defparam GSB_CNT_3_48_0_inst.sps_h6w6.CONF = "101";
  defparam GSB_CNT_3_48_0_inst.sps_h6w8.CONF = "101";
  defparam GSB_CNT_3_48_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_48_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_48_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_48_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_48_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_48_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_48_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_48_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_48_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(\net_Buf-pad-RGB[23]_RIGHT_H6W4_to_H6E43_48_0 ),
    .H6E5(),
    .H6E6(\net_Buf-pad-RGB[20]_RIGHT_H6W6_to_H6E63_48_0 ),
    .H6E7(),
    .H6E8(\net_Buf-pad-RGB[23]_RIGHT_H6W8_to_H6E83_48_0 ),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(\net_Buf-pad-RGB[23]_H6W4_to_H6E43_42_0 ),
    .H6W5(),
    .H6W6(\net_Buf-pad-RGB[20]_H6W6_to_H6E63_42_0 ),
    .H6W7(),
    .H6W8(\net_Buf-pad-RGB[23]_H6W8_to_H6E83_42_0 ),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_40_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_40_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_40_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6e0.CONF = "01011011";
  defparam GSB_TOP_1_40_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s16.CONF = "01";
  defparam GSB_TOP_1_40_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6s6.CONF = "111011";
  defparam GSB_TOP_1_40_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_40_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_40_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6a3.CONF = "01011";
  defparam GSB_TOP_1_40_0_inst.sps_v6b0.CONF = "01101";
  defparam GSB_TOP_1_40_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d0.CONF = "01101";
  defparam GSB_TOP_1_40_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d10.CONF = "110111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_40_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_40_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_40_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(\net_Buf-pad-RGB[6]_TOP_S16_to_N162_40_0 ),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(\net_Buf-pad-RGB[12]_TOP_H6E0_to_TOP_H6M01_44_0 ),
    .TOP_H6E1(\net_Buf-pad-RGB[4]_TOP_H6W1_to_TOP_H6E11_40_0 ),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(\net_Buf-pad-RGB[6]_TOP_H6W2_to_TOP_H6M21_40_0 ),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(\net_Buf-pad-RGB[13]_TOP_V6A3_to_V6N32_40_0 ),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(\net_Buf-pad-RGB[13]_TOP_V6B0_to_V6N03_40_0 ),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(\net_Buf-pad-RGB[12]_TOP_V6D0_to_V6M03_40_0 ),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(\net_Buf-pad-RGB[6]_TOP_V6D10_to_V6M103_40_0 ),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(\net_Buf-pad-RGB[4]_TOP_V6S6_to_V6M64_40_0 ),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(\net_Buf-pad-RGB[13]_IN_to_TOP_I21_40_0 ),
    .TOP_I1(\net_Buf-pad-RGB[12]_IN_to_TOP_I11_40_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_CNT_2_40_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_2_40_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_2_40_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_s22.CONF = "01";
  defparam GSB_CNT_2_40_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_2_40_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_2_40_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_2_40_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_2_40_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s16_n16.CONF = "0";
  defparam GSB_CNT_2_40_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s21_e23.CONF = "0";
  defparam GSB_CNT_2_40_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s9_e11.CONF = "0";
  defparam GSB_CNT_2_40_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_2_40_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_2_40_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(\net_Buf-pad-RGB[22]_W11_to_E112_40_0 ),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(\net_Buf-pad-RGB[22]_W23_to_E232_40_0 ),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(\net_Buf-pad-RGB[6]_TOP_S16_to_N162_40_0 ),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(\net_Buf-pad-RGB[22]_S9_to_N93_40_0 ),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(\net_Buf-pad-RGB[6]_S16_to_N163_40_0 ),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(\net_Buf-pad-RGB[22]_S21_to_N213_40_0 ),
    .S22(\net_Buf-pad-RGB[13]_S22_to_N223_40_0 ),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(\net_Buf-pad-RGB[13]_TOP_V6A3_to_V6N32_40_0 ),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_50_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w2.CONF = "01011011";
  defparam GSB_TOP_1_50_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_50_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_50_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_50_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_50_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_50_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_50_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_50_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(\net_Buf-pad-RGB[6]_TOP_H6W2_to_TOP_H6E21_44_0 ),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(\net_Buf-pad-RGB[6]_IN_to_TOP_I11_50_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_44_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w1.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w2.CONF = "01101110";
  defparam GSB_TOP_1_44_0_inst.sps_h6w3.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w4.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_44_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_44_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s2.CONF = "0101111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_44_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_44_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d6.CONF = "110111";
  defparam GSB_TOP_1_44_0_inst.sps_v6d8.CONF = "110111";
  defparam GSB_TOP_1_44_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_44_0_inst.sps_v6m1.CONF = "01101";
  defparam GSB_TOP_1_44_0_inst.sps_v6m2.CONF = "01110";
  defparam GSB_TOP_1_44_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_44_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(\net_Buf-pad-RGB[6]_TOP_H6W2_to_TOP_H6E21_44_0 ),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(\net_Buf-pad-RGB[12]_TOP_H6E0_to_TOP_H6M01_44_0 ),
    .TOP_H6M1(\net_Buf-pad-RGB[4]_TOP_H6W1_to_TOP_H6E11_40_0 ),
    .TOP_H6M2(),
    .TOP_H6M3(\net_Buf-pad-RGB[5]_TOP_H6W3_to_TOP_H6M31_44_0 ),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(),
    .TOP_H6W2(\net_Buf-pad-RGB[6]_TOP_H6W2_to_TOP_H6M21_40_0 ),
    .TOP_H6W3(),
    .TOP_H6W4(),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(\net_Buf-pad-RGB[10]_TOP_V6M1_to_V6N14_44_0 ),
    .TOP_V6M2(\net_Buf-pad-RGB[10]_TOP_V6M2_to_V6N24_44_0 ),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(\net_Buf-pad-RGB[12]_TOP_V6D6_to_V6M63_44_0 ),
    .TOP_V6D7(),
    .TOP_V6D8(\net_Buf-pad-RGB[5]_TOP_V6D8_to_V6M83_44_0 ),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(\net_Buf-pad-RGB[4]_TOP_V6S2_to_V6M24_44_0 ),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(),
    .TOP_I1(\net_Buf-pad-RGB[10]_IN_to_TOP_I11_44_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_RHT_30_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_30_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_30_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_30_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_30_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_30_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_30_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_30_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_llv0.CONF = "0011011111";
  defparam GSB_RHT_30_54_0_inst.sps_llv6.CONF = "0001111111";
  defparam GSB_RHT_30_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_30_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_30_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_30_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_30_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_30_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_30_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_30_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_30_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_30_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_30_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_30_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_30_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_30_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_30_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_30_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_30_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(\net_Buf-pad-RGB[21]_RIGHT_LLV0_to_RIGHT_LLV05_54_0 ),
    .RIGHT_LLV6(\net_Buf-pad-RGB[22]_RIGHT_LLV6_to_RIGHT_LLV65_54_0 ),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(\net_Buf-pad-RGB[21]_IN_to_RIGHT_I230_54_0 ),
    .RIGHT_I3(\net_Buf-pad-RGB[22]_IN_to_RIGHT_I330_54_0 ),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_RHT_2_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_2_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_2_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_2_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_2_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_2_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_2_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_2_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_2_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6d4.CONF = "110111";
  defparam GSB_RHT_2_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_2_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_2_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_2_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_h6w10.CONF = "110111";
  defparam GSB_RHT_2_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_2_54_0_inst.sps_h6w6.CONF = "110111";
  defparam GSB_RHT_2_54_0_inst.sps_h6w8.CONF = "110111";
  defparam GSB_RHT_2_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_2_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_2_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_2_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_2_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_2_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_2_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_2_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_2_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_2_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_2_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_2_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_2_54_0_inst.sps_v6s0.CONF = "00111011";
  defparam GSB_RHT_2_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_2_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_2_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_2_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_2_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_2_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_2_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_2_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_2_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_2_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_2_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_2_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_2_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(\net_Buf-pad-RGB[21]_RIGHT_H6D4_to_H6E42_49_0 ),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(\net_Buf-pad-RGB[21]_RIGHT_H6W6_to_H6E62_48_0 ),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(\net_Buf-pad-RGB[22]_RIGHT_H6W8_to_H6E82_48_0 ),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(\net_Buf-pad-RGB[22]_RIGHT_H6W10_to_H6E102_48_0 ),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(\net_Buf-pad-RGB[21]_RIGHT_V6N0_to_RIGHT_V6M02_54_0 ),
    .RIGHT_V6M1(\net_Buf-pad-RGB[21]_RIGHT_V6N1_to_RIGHT_V6M12_54_0 ),
    .RIGHT_V6M2(\net_Buf-pad-RGB[22]_RIGHT_V6N2_to_RIGHT_V6M22_54_0 ),
    .RIGHT_V6M3(\net_Buf-pad-RGB[22]_RIGHT_V6N3_to_RIGHT_V6M32_54_0 ),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(\net_Buf-pad-RGB[18]_RIGHT_V6S0_to_RIGHT_V6M05_54_0 ),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(\net_Buf-pad-RGB[18]_RIGHT_LLV0_to_RIGHT_LLV02_54_0 ),
    .RIGHT_LLV6(),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(),
    .RIGHT_I3(),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_2_48_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_h6w10.CONF = "101";
  defparam GSB_CNT_2_48_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_h6w6.CONF = "101";
  defparam GSB_CNT_2_48_0_inst.sps_h6w8.CONF = "101";
  defparam GSB_CNT_2_48_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_2_48_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_2_48_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_2_48_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_2_48_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_2_48_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_2_48_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_2_48_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_2_48_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(\net_Buf-pad-RGB[21]_RIGHT_H6W6_to_H6E62_48_0 ),
    .H6E7(),
    .H6E8(\net_Buf-pad-RGB[22]_RIGHT_H6W8_to_H6E82_48_0 ),
    .H6E9(),
    .H6E10(\net_Buf-pad-RGB[22]_RIGHT_H6W10_to_H6E102_48_0 ),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_Buf-pad-RGB[21]_H6W6_to_H6E62_42_0 ),
    .H6W7(),
    .H6W8(\net_Buf-pad-RGB[22]_H6W8_to_H6E82_42_0 ),
    .H6W9(),
    .H6W10(\net_Buf-pad-RGB[22]_H6W10_to_H6E102_42_0 ),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_2_42_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_2_42_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_2_42_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_v6n0.CONF = "0010";
  defparam GSB_CNT_2_42_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w11.CONF = "01";
  defparam GSB_CNT_2_42_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w23.CONF = "01";
  defparam GSB_CNT_2_42_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s15.CONF = "01";
  defparam GSB_CNT_2_42_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_s2.CONF = "01";
  defparam GSB_CNT_2_42_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_2_42_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_2_42_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_2_42_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_2_42_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_2_42_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_2_42_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(\net_Buf-pad-RGB[22]_W11_to_E112_40_0 ),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(\net_Buf-pad-RGB[22]_W23_to_E232_40_0 ),
    .S0(),
    .S1(),
    .S2(\net_Buf-pad-RGB[5]_S2_to_N23_42_0 ),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(\net_Buf-pad-RGB[21]_S15_to_N153_42_0 ),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(\net_Buf-pad-RGB[21]_H6W6_to_H6E62_42_0 ),
    .H6E7(),
    .H6E8(\net_Buf-pad-RGB[22]_H6W8_to_H6E82_42_0 ),
    .H6E9(),
    .H6E10(\net_Buf-pad-RGB[22]_H6W10_to_H6E102_42_0 ),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(\net_Buf-pad-RGB[5]_TOP_LLV11_to_LLV02_42_0 ),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_3_44_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_44_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_44_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_w13.CONF = "0";
  defparam GSB_CNT_3_44_0_inst.sps_w14.CONF = "0";
  defparam GSB_CNT_3_44_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_44_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_44_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_44_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_44_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_44_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_44_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(\net_Buf-pad-RGB[5]_W13_to_E133_43_0 ),
    .W14(\net_Buf-pad-RGB[12]_W14_to_E143_43_0 ),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(\net_Buf-pad-RGB[12]_TOP_V6D6_to_V6M63_44_0 ),
    .V6M7(),
    .V6M8(\net_Buf-pad-RGB[5]_TOP_V6D8_to_V6M83_44_0 ),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_3_43_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_43_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_43_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w11.CONF = "10";
  defparam GSB_CNT_3_43_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_out2.CONF = "000111";
  defparam GSB_CNT_3_43_0_inst.sps_out3.CONF = "000111";
  defparam GSB_CNT_3_43_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_s0_bx_b.CONF = "001011";
  defparam GSB_CNT_3_43_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s0_f_b1.CONF = "010111101";
  defparam GSB_CNT_3_43_0_inst.sps_s0_f_b2.CONF = "100011111";
  defparam GSB_CNT_3_43_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_43_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_43_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_s3.CONF = "01";
  defparam GSB_CNT_3_43_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s7.CONF = "0";
  defparam GSB_CNT_3_43_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_43_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_43_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_43_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_43_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n3_w4.CONF = "0";
  defparam GSB_CNT_3_43_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_43_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_43_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(\net_Buf-pad-RGB[5]_W13_to_E133_43_0 ),
    .E14(\net_Buf-pad-RGB[12]_W14_to_E143_43_0 ),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(\net_Buf-pad-RGB[21]_S3_to_N33_43_0 ),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(net_U18_S_W11_to_E113_42_0),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(\net_Buf-pad-RGB[20]_S3_to_N34_43_0 ),
    .S4(),
    .S5(),
    .S6(),
    .S7(net_U18_S_S7_to_N74_43_0),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(\net_Buf-pad-RGB[20]_H6W4_to_H6E43_43_0 ),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-RGB[12]_S0_F_B1_to_F13_43_0 ),
    .S0_F_B2(\net_Buf-pad-RGB[5]_S0_F_B2_to_F23_43_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(\net_Buf-pad-RGB[21]_S0_BX_B_to_BX3_43_0 ),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(net_U18_S_X_to_S0_X3_43_0),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_TOP_1_53_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6w1.CONF = "01011011";
  defparam GSB_TOP_1_53_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6w3.CONF = "01011110";
  defparam GSB_TOP_1_53_0_inst.sps_h6w4.CONF = "01101011";
  defparam GSB_TOP_1_53_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_53_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_53_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6s8.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_53_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_53_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6c2.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_53_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_53_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_53_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(),
    .TOP_H6E2(),
    .TOP_H6E3(),
    .TOP_H6E4(),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(\net_Buf-pad-RGB[4]_TOP_H6W1_to_TOP_H6E11_47_0 ),
    .TOP_H6W2(),
    .TOP_H6W3(\net_Buf-pad-RGB[5]_TOP_H6W3_to_TOP_H6E31_47_0 ),
    .TOP_H6W4(\net_Buf-pad-RGB[5]_TOP_H6W4_to_TOP_H6E41_47_0 ),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(\net_Buf-pad-RGB[5]_IN_to_TOP_I21_53_0 ),
    .TOP_I1(\net_Buf-pad-RGB[4]_IN_to_TOP_I11_53_0 ),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_TOP_1_47_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6w0.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6w1.CONF = "01101110";
  defparam GSB_TOP_1_47_0_inst.sps_h6w2.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6w3.CONF = "01101110";
  defparam GSB_TOP_1_47_0_inst.sps_h6w4.CONF = "01110110";
  defparam GSB_TOP_1_47_0_inst.sps_ice1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_ice2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_llh0.CONF = "1111111111";
  defparam GSB_TOP_1_47_0_inst.sps_llh6.CONF = "1111111111";
  defparam GSB_TOP_1_47_0_inst.sps_llv0.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv6.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_o1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_o2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_oce1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_oce2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_sr_b1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_sr_b2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_t1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_t2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_tce1.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_tce2.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s0.CONF = "1111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s1.CONF = "1111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s2.CONF = "1111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s3.CONF = "1111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e0.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e1.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e2.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e3.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6e5.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_s0.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s1.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s10.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s11.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s12.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s13.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s14.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s15.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s16.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s17.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s18.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s19.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s2.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s20.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s21.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s22.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s23.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s3.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s4.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s5.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s6.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s7.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s8.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_s9.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_v6s10.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s4.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s6.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6s8.CONF = "111101";
  defparam GSB_TOP_1_47_0_inst.sps_llv4.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv8.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv1.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv5.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv9.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_h6e4.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_h6w5.CONF = "11111111";
  defparam GSB_TOP_1_47_0_inst.sps_llv10.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv11.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv2.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv3.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_llv7.CONF = "11";
  defparam GSB_TOP_1_47_0_inst.sps_v6a0.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6a1.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6a2.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6a3.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6b0.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6b1.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6b2.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6b3.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6c0.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6c1.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6c2.CONF = "01101";
  defparam GSB_TOP_1_47_0_inst.sps_v6c3.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d0.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d1.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d10.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d2.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d3.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d4.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d6.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6d8.CONF = "111111";
  defparam GSB_TOP_1_47_0_inst.sps_v6m0.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6m1.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6m2.CONF = "11111";
  defparam GSB_TOP_1_47_0_inst.sps_v6m3.CONF = "11111";
  GSB_TOP GSB_TOP_1_47_0_inst (
    .TOP_S23(),
    .TOP_S22(),
    .TOP_S21(),
    .TOP_S20(),
    .TOP_S19(),
    .TOP_S18(),
    .TOP_S17(),
    .TOP_S16(),
    .TOP_S15(),
    .TOP_S14(),
    .TOP_S13(),
    .TOP_S12(),
    .TOP_S11(),
    .TOP_S10(),
    .TOP_S9(),
    .TOP_S8(),
    .TOP_S7(),
    .TOP_S6(),
    .TOP_S5(),
    .TOP_S4(),
    .TOP_S3(),
    .TOP_S2(),
    .TOP_S1(),
    .TOP_S0(),
    .TOP_H6E0(),
    .TOP_H6E1(\net_Buf-pad-RGB[4]_TOP_H6W1_to_TOP_H6E11_47_0 ),
    .TOP_H6E2(),
    .TOP_H6E3(\net_Buf-pad-RGB[5]_TOP_H6W3_to_TOP_H6E31_47_0 ),
    .TOP_H6E4(\net_Buf-pad-RGB[5]_TOP_H6W4_to_TOP_H6E41_47_0 ),
    .TOP_H6E5(),
    .TOP_H6A0(),
    .TOP_H6A1(),
    .TOP_H6A2(),
    .TOP_H6A3(),
    .TOP_H6A4(),
    .TOP_H6A5(),
    .TOP_H6B0(),
    .TOP_H6B1(),
    .TOP_H6B2(),
    .TOP_H6B3(),
    .TOP_H6B4(),
    .TOP_H6B5(),
    .TOP_H6M0(),
    .TOP_H6M1(),
    .TOP_H6M2(),
    .TOP_H6M3(),
    .TOP_H6M4(),
    .TOP_H6M5(),
    .TOP_H6C0(),
    .TOP_H6C1(),
    .TOP_H6C2(),
    .TOP_H6C3(),
    .TOP_H6C4(),
    .TOP_H6C5(),
    .TOP_H6D0(),
    .TOP_H6D1(),
    .TOP_H6D2(),
    .TOP_H6D3(),
    .TOP_H6D4(),
    .TOP_H6D5(),
    .TOP_H6W0(),
    .TOP_H6W1(\net_Buf-pad-RGB[4]_TOP_H6W1_to_TOP_H6E11_40_0 ),
    .TOP_H6W2(),
    .TOP_H6W3(\net_Buf-pad-RGB[5]_TOP_H6W3_to_TOP_H6M31_44_0 ),
    .TOP_H6W4(\net_Buf-pad-RGB[5]_TOP_H6W4_to_TOP_H6A41_42_0 ),
    .TOP_H6W5(),
    .TOP_V6A0(),
    .TOP_V6A1(),
    .TOP_V6A2(),
    .TOP_V6A3(),
    .TOP_V6A4(),
    .TOP_V6A5(),
    .TOP_V6A6(),
    .TOP_V6A7(),
    .TOP_V6A8(),
    .TOP_V6A9(),
    .TOP_V6A10(),
    .TOP_V6A11(),
    .TOP_V6B0(),
    .TOP_V6B1(),
    .TOP_V6B2(),
    .TOP_V6B3(),
    .TOP_V6B4(),
    .TOP_V6B5(),
    .TOP_V6B6(),
    .TOP_V6B7(),
    .TOP_V6B8(),
    .TOP_V6B9(),
    .TOP_V6B10(),
    .TOP_V6B11(),
    .TOP_V6M0(),
    .TOP_V6M1(),
    .TOP_V6M2(),
    .TOP_V6M3(),
    .TOP_V6M4(),
    .TOP_V6M5(),
    .TOP_V6M6(),
    .TOP_V6M7(),
    .TOP_V6M8(),
    .TOP_V6M9(),
    .TOP_V6M10(),
    .TOP_V6M11(),
    .TOP_V6C0(),
    .TOP_V6C1(),
    .TOP_V6C2(\net_Buf-pad-RGB[9]_TOP_V6C2_to_V6N25_47_0 ),
    .TOP_V6C3(),
    .TOP_V6C4(),
    .TOP_V6C5(),
    .TOP_V6C6(),
    .TOP_V6C7(),
    .TOP_V6C8(),
    .TOP_V6C9(),
    .TOP_V6C10(),
    .TOP_V6C11(),
    .TOP_V6D0(),
    .TOP_V6D1(),
    .TOP_V6D2(),
    .TOP_V6D3(),
    .TOP_V6D4(),
    .TOP_V6D5(),
    .TOP_V6D6(),
    .TOP_V6D7(),
    .TOP_V6D8(),
    .TOP_V6D9(),
    .TOP_V6D10(),
    .TOP_V6D11(),
    .TOP_V6S0(),
    .TOP_V6S1(),
    .TOP_V6S2(),
    .TOP_V6S3(),
    .TOP_V6S4(),
    .TOP_V6S5(),
    .TOP_V6S6(),
    .TOP_V6S7(),
    .TOP_V6S8(\net_Buf-pad-RGB[9]_TOP_V6S8_to_V6M84_47_0 ),
    .TOP_V6S9(),
    .TOP_V6S10(),
    .TOP_V6S11(),
    .TOP_LLH0(),
    .TOP_LLH6(),
    .TOP_LLV0(),
    .TOP_LLV1(),
    .TOP_LLV2(),
    .TOP_LLV3(),
    .TOP_LLV4(),
    .TOP_LLV5(),
    .TOP_LLV6(),
    .TOP_LLV7(),
    .TOP_LLV8(),
    .TOP_LLV9(),
    .TOP_LLV10(),
    .TOP_LLV11(),
    .TOP_HGCLK0(),
    .TOP_HGCLK1(),
    .TOP_HGCLK2(),
    .TOP_HGCLK3(),
    .TOP_I2(\net_Buf-pad-RGB[9]_IN_to_TOP_I21_47_0 ),
    .TOP_I1(),
    .TOP_IQ2(),
    .TOP_IQ1(),
    .TOP_ICE2(),
    .TOP_ICE1(),
    .TOP_O2(),
    .TOP_O1(),
    .TOP_OCE2(),
    .TOP_OCE1(),
    .TOP_T2(),
    .TOP_T1(),
    .TOP_TCE2(),
    .TOP_TCE1(),
    .TOP_CLK2(),
    .TOP_CLK1(),
    .TOP_SR_B2(),
    .TOP_SR_B1()
  );

  defparam GSB_CNT_2_49_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_h6w4.CONF = "101";
  defparam GSB_CNT_2_49_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_2_49_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_2_49_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_2_49_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_2_49_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_2_49_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_2_49_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_2_49_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_2_49_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(\net_Buf-pad-RGB[21]_RIGHT_H6D4_to_H6E42_49_0 ),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(\net_Buf-pad-RGB[21]_H6W4_to_H6E42_43_0 ),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_2_43_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_2_43_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_2_43_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_s3.CONF = "01";
  defparam GSB_CNT_2_43_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_2_43_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_2_43_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_2_43_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_2_43_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_2_43_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_2_43_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(\net_Buf-pad-RGB[21]_S3_to_N33_43_0 ),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(\net_Buf-pad-RGB[21]_H6W4_to_H6E42_43_0 ),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_43_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_43_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_43_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_w10.CONF = "10";
  defparam GSB_CNT_4_43_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_out1.CONF = "000111";
  defparam GSB_CNT_4_43_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_out3.CONF = "000111";
  defparam GSB_CNT_4_43_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_s0_bx_b.CONF = "001011";
  defparam GSB_CNT_4_43_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s0_f_b1.CONF = "001111011";
  defparam GSB_CNT_4_43_0_inst.sps_s0_f_b2.CONF = "001011111";
  defparam GSB_CNT_4_43_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_43_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_43_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_43_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_43_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_43_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_43_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e11_w11.CONF = "0";
  defparam GSB_CNT_4_43_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n3_w4.CONF = "0";
  defparam GSB_CNT_4_43_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n7_w8.CONF = "0";
  defparam GSB_CNT_4_43_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_43_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_43_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(\net_Lut-U21_0_0_W11_to_E114_43_0 ),
    .E12(),
    .E13(),
    .E14(),
    .E15(\net_Buf-pad-RGB[4]_W15_to_E154_43_0 ),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(\net_Buf-pad-RGB[20]_S3_to_N34_43_0 ),
    .N4(),
    .N5(),
    .N6(),
    .N7(net_U18_S_S7_to_N74_43_0),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(\net_Buf-pad-RGB[11]_E7_to_W74_43_0 ),
    .W8(net_U18_S_W8_to_E84_42_0),
    .W9(),
    .W10(net_U23_S_W10_to_E104_42_0),
    .W11(\net_Lut-U21_0_0_W11_to_E114_42_0 ),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(net_U23_S_OUT1_to_OUT_W14_44_0),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Buf-pad-RGB[11]_S0_F_B1_to_F14_43_0 ),
    .S0_F_B2(\net_Buf-pad-RGB[4]_S0_F_B2_to_F24_43_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(\net_Buf-pad-RGB[20]_S0_BX_B_to_BX4_43_0 ),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(net_U23_S_X_to_S0_X4_43_0),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_40_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_40_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_40_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e12.CONF = "10";
  defparam GSB_CNT_4_40_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_40_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_40_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_40_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_40_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s10_e4.CONF = "0";
  defparam GSB_CNT_4_40_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_40_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_40_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(net_U20_CO_E4_to_W44_42_0),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(\net_Buf-pad-RGB[4]_E12_to_W124_42_0 ),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(net_U20_CO_N10_to_S104_40_0),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(\net_Buf-pad-RGB[4]_TOP_V6S6_to_V6M64_40_0 ),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_RHT_28_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_28_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_28_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_28_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_28_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_28_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_28_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_28_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_28_54_0_inst.sps_llv6.CONF = "0001111111";
  defparam GSB_RHT_28_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_28_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_28_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_28_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_28_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_28_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_28_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_28_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_28_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_28_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_28_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_28_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_28_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_28_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_28_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_28_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_28_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(),
    .RIGHT_LLV6(\net_Buf-pad-RGB[20]_RIGHT_LLV6_to_UR_LLV41_54_0 ),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(),
    .RIGHT_I3(\net_Buf-pad-RGB[20]_IN_to_RIGHT_I328_54_0 ),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_UR_1_54_0_inst.sps_h6a0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6a1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6a2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6a3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6b0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6b1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6b2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6b3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6c0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6c1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6c2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6c3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6d0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6d1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6d2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6d3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6d4.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6m0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6m1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6m2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6m3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6w0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6w1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6w2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6w3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6w4.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_llv0.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_llv6.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_v6s0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6s1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6s2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6s3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6a5.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_llv4.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_llv8.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_llv1.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_llv5.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_llv9.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_h6w5.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_llv10.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_llv11.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_llv2.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_llv3.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_llv7.CONF = "1";
  defparam GSB_UR_1_54_0_inst.sps_v6a0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6a1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6a2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6a3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6b0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6b1.CONF = "00";
  defparam GSB_UR_1_54_0_inst.sps_v6b2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6b3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6c0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6c1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6c2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6c3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6d0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6d1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6d2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6d3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6m0.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6m1.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6m2.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_v6m3.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6a4.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6b4.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6b5.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6c4.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6c5.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6d5.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6m4.CONF = "11";
  defparam GSB_UR_1_54_0_inst.sps_h6m5.CONF = "11";
  GSB_UR GSB_UR_1_54_0_inst (
    .UR_H6W0(),
    .UR_H6D0(),
    .UR_H6C0(),
    .UR_H6M0(),
    .UR_H6B0(),
    .UR_H6A0(),
    .UR_H6W1(),
    .UR_H6D1(),
    .UR_H6C1(),
    .UR_H6M1(),
    .UR_H6B1(),
    .UR_H6A1(),
    .UR_H6W2(),
    .UR_H6D2(),
    .UR_H6C2(),
    .UR_H6M2(),
    .UR_H6B2(),
    .UR_H6A2(),
    .UR_H6W3(),
    .UR_H6D3(),
    .UR_H6C3(),
    .UR_H6M3(),
    .UR_H6B3(),
    .UR_H6A3(),
    .UR_H6W4(),
    .UR_H6D4(),
    .UR_H6C4(),
    .UR_H6M4(),
    .UR_H6B4(),
    .UR_H6A4(),
    .UR_H6W5(),
    .UR_H6D5(),
    .UR_H6C5(),
    .UR_H6M5(),
    .UR_H6B5(),
    .UR_H6A5(),
    .UR_LLH0(),
    .UR_LLH1(),
    .UR_LLH2(),
    .UR_LLH3(),
    .UR_LLH4(),
    .UR_LLH5(),
    .UR_LLH6(),
    .UR_LLH7(),
    .UR_LLH8(),
    .UR_LLH9(),
    .UR_LLH10(),
    .UR_LLH11(),
    .UR_V6S0(),
    .UR_V6D0(),
    .UR_V6C0(),
    .UR_V6M0(),
    .UR_V6B0(),
    .UR_V6A0(),
    .UR_V6S1(),
    .UR_V6D1(),
    .UR_V6C1(),
    .UR_V6M1(),
    .UR_V6B1(\net_Buf-pad-RGB[20]_UR_V6B1_to_RIGHT_V6N13_54_0 ),
    .UR_V6A1(),
    .UR_V6S2(),
    .UR_V6D2(),
    .UR_V6C2(),
    .UR_V6M2(),
    .UR_V6B2(),
    .UR_V6A2(),
    .UR_V6S3(),
    .UR_V6D3(),
    .UR_V6C3(),
    .UR_V6M3(),
    .UR_V6B3(),
    .UR_V6A3(),
    .UR_LLV0(),
    .UR_LLV1(),
    .UR_LLV2(),
    .UR_LLV3(),
    .UR_LLV4(\net_Buf-pad-RGB[20]_RIGHT_LLV6_to_UR_LLV41_54_0 ),
    .UR_LLV5(),
    .UR_LLV6(),
    .UR_LLV7(),
    .UR_LLV8(),
    .UR_LLV9(),
    .UR_LLV10(),
    .UR_LLV11()
  );

  defparam GSB_CNT_3_49_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_h6w4.CONF = "101";
  defparam GSB_CNT_3_49_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_3_49_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_3_49_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_3_49_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_3_49_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_3_49_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_3_49_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_3_49_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_3_49_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(\net_Buf-pad-RGB[20]_RIGHT_H6D4_to_H6E43_49_0 ),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(\net_Buf-pad-RGB[20]_H6W4_to_H6E43_43_0 ),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_40_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_40_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_40_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n10.CONF = "10";
  defparam GSB_CNT_5_40_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_40_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_40_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_40_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_40_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_40_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_40_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(net_U20_CO_N10_to_S104_40_0),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(net_U20_CO_H6W1_to_H6M15_40_0),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_49_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_h6w6.CONF = "101";
  defparam GSB_CNT_5_49_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_49_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_49_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_49_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_49_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_49_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_49_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_49_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_49_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(\net_Buf-pad-RGB[18]_RIGHT_H6D6_to_H6E65_49_0 ),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_Buf-pad-RGB[18]_H6W6_to_H6E65_43_0 ),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_43_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_43_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_43_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s15.CONF = "01";
  defparam GSB_CNT_5_43_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_43_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_43_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_43_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_43_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s15_e13.CONF = "0";
  defparam GSB_CNT_5_43_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_43_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_43_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(\net_Buf-pad-RGB[18]_E13_to_W135_44_0 ),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(\net_Buf-pad-RGB[18]_H6W6_to_H6E65_43_0 ),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_48_0_inst.sps_h6w0.CONF = "0000";
  defparam GSB_CNT_5_48_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_48_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_48_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_48_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_48_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_48_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_48_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_48_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_48_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(\net_Buf-pad-RGB[18]_RIGHT_H6W0_to_H6E05_48_0 ),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(\net_Buf-pad-RGB[18]_H6W0_to_H6M05_45_0 ),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_RHT_6_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_6_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_6_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_6_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_6_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6c2.CONF = "01110";
  defparam GSB_RHT_6_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6d8.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w0.CONF = "0111101";
  defparam GSB_RHT_6_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_6_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh2.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh3.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_6_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_6_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_6_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_6_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_6_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_6_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_6_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_6_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_6_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_6_54_0_inst.sps_w9.CONF = "111";
  GSB_RHT GSB_RHT_6_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(\net_Buf-pad-RGB[2]_RIGHT_H6C2_to_H6E26_50_0 ),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(\net_Buf-pad-RGB[2]_RIGHT_H6W0_to_H6E06_48_0 ),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(),
    .RIGHT_LLH3(),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(),
    .RIGHT_LLV6(),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(\net_Buf-pad-RGB[2]_IN_to_RIGHT_I16_54_0 ),
    .RIGHT_I2(),
    .RIGHT_I3(),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_6_50_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_h6w2.CONF = "0000";
  defparam GSB_CNT_6_50_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_50_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_50_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_50_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_50_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_50_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_50_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_50_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_50_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(\net_Buf-pad-RGB[2]_RIGHT_H6C2_to_H6E26_50_0 ),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(\net_Buf-pad-RGB[2]_H6W2_to_H6E26_44_0 ),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_44_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_44_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_44_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_v6s3.CONF = "0100";
  defparam GSB_CNT_6_44_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n19.CONF = "01";
  defparam GSB_CNT_6_44_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_44_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_44_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_44_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_44_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_44_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_44_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(\net_Buf-pad-RGB[2]_N19_to_S195_44_0 ),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(\net_Buf-pad-RGB[2]_H6W2_to_H6E26_44_0 ),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_48_0_inst.sps_h6w0.CONF = "0000";
  defparam GSB_CNT_6_48_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_48_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_48_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_48_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_48_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_48_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_48_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_48_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_48_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(\net_Buf-pad-RGB[2]_RIGHT_H6W0_to_H6E06_48_0 ),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(\net_Buf-pad-RGB[2]_H6W0_to_H6M06_45_0 ),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_45_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_45_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_45_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_n4.CONF = "10";
  defparam GSB_CNT_6_45_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_45_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_45_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_45_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_45_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_45_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_45_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(\net_Buf-pad-RGB[2]_N4_to_S45_45_0 ),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(\net_Buf-pad-RGB[2]_H6W0_to_H6M06_45_0 ),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_46_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_46_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_46_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_46_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_46_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_46_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_46_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n20_e16.CONF = "0";
  defparam GSB_CNT_5_46_0_inst.switch_n20_w1.CONF = "0";
  defparam GSB_CNT_5_46_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_46_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_46_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(\net_Buf-pad-RGB[9]_W16_to_E165_46_0 ),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(\net_Buf-pad-RGB[9]_W1_to_E15_45_0 ),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );
endmodule
