
module display (clk, rst_n, lcd_db, lcd_en, lcd_rs, lcd_rw, lcd_rst);
 input clk;
 input rst_n;
 output [7:0] lcd_db;
 output lcd_en;
 output lcd_rs;
 output lcd_rw;
 output lcd_rst;
  wire \net_cnt_lcd_reg[6]_XQ_to_S1_XQ7_6_0 ;
  wire \net_cnt_lcd_reg[6]_H6E7_to_H6M77_9_0 ;
  wire \net_cnt_lcd_reg[6]_S1_G_B3_to_G37_9_0 ;
  wire \net_cnt_lcd_reg[6]_E14_to_W147_7_0 ;
  wire \net_cnt_lcd_reg[6]_E14_to_W147_8_0 ;
  wire \net_cnt_lcd_reg[6]_S0_F_B4_to_F47_8_0 ;
  wire \net_cnt_lcd_reg[6]_S13_to_N138_6_0 ;
  wire \net_cnt_lcd_reg[6]_E13_to_W138_7_0 ;
  wire \net_cnt_lcd_reg[6]_S0_F_B4_to_F48_7_0 ;
  wire \net_cnt_lcd_reg[6]_S17_to_N178_9_0 ;
  wire \net_cnt_lcd_reg[6]_S0_F_B3_to_F38_9_0 ;
  wire \net_cnt_lcd_reg[6]_E17_to_W177_10_0 ;
  wire \net_cnt_lcd_reg[6]_S1_F_B3_to_F37_10_0 ;
  wire \net_cnt_lcd_reg[6]_V6S6_to_V6M610_9_0 ;
  wire \net_cnt_lcd_reg[6]_E12_to_W1210_10_0 ;
  wire \net_cnt_lcd_reg[6]_S0_G_B3_to_G310_10_0 ;
  wire \net_cnt_lcd_reg[6]_H6E3_to_H6M37_9_0 ;
  wire \net_cnt_lcd_reg[6]_S0_F_B3_to_F37_9_0 ;
  wire \net_cnt_lcd_reg[6]_S1_F_B2_to_F210_10_0 ;
  wire \net_cnt_lcd_reg[6]_S17_to_N179_9_0 ;
  wire \net_cnt_lcd_reg[6]_S0_G_B2_to_G29_9_0 ;
  wire \net_cnt_lcd_reg[6]_S1_G_B3_to_G38_7_0 ;
  wire \net_cnt_lcd_reg[6]_V6S2_to_V6M210_6_0 ;
  wire \net_cnt_lcd_reg[6]_H6E2_to_H6M210_9_0 ;
  wire \net_cnt_lcd_reg[6]_S0_F_B2_to_F210_9_0 ;
  wire \net_cnt_lcd_reg[6]_S0_G_B2_to_G210_9_0 ;
  wire \net_cnt_lcd_reg[6]_W19_to_E197_5_0 ;
  wire \net_cnt_lcd_reg[6]_S0_F_B1_to_F17_5_0 ;
  wire \net_cnt_lcd_reg[0]_XQ_to_S1_XQ7_5_0 ;
  wire \net_cnt_lcd_reg[0]_H6E3_to_H6M37_8_0 ;
  wire \net_cnt_lcd_reg[0]_E21_to_W217_9_0 ;
  wire \net_cnt_lcd_reg[0]_S1_G_B4_to_G47_9_0 ;
  wire \net_cnt_lcd_reg[0]_S22_to_N228_5_0 ;
  wire \net_cnt_lcd_reg[0]_E18_to_W188_6_0 ;
  wire \net_cnt_lcd_reg[0]_S16_to_N169_6_0 ;
  wire \net_cnt_lcd_reg[0]_S0_G_B2_to_G29_6_0 ;
  wire \net_cnt_lcd_reg[0]_H6E5_to_H6M57_8_0 ;
  wire \net_cnt_lcd_reg[0]_S4_to_N48_8_0 ;
  wire \net_cnt_lcd_reg[0]_E0_to_W08_9_0 ;
  wire \net_cnt_lcd_reg[0]_S0_F_B4_to_F48_9_0 ;
  wire \net_cnt_lcd_reg[0]_W20_to_E207_10_0 ;
  wire \net_cnt_lcd_reg[0]_S1_F_B4_to_F47_10_0 ;
  wire \net_cnt_lcd_reg[0]_V6S3_to_V6M310_11_0 ;
  wire \net_cnt_lcd_reg[0]_W20_to_E2010_10_0 ;
  wire \net_cnt_lcd_reg[0]_S0_G_B4_to_G410_10_0 ;
  wire \net_cnt_lcd_reg[0]_E2_to_W27_9_0 ;
  wire \net_cnt_lcd_reg[0]_S0_F_B4_to_F47_9_0 ;
  wire \net_cnt_lcd_reg[0]_W18_to_E1810_10_0 ;
  wire \net_cnt_lcd_reg[0]_S1_F_B3_to_F310_10_0 ;
  wire \net_cnt_lcd_reg[0]_V6S3_to_V6M310_8_0 ;
  wire \net_cnt_lcd_reg[0]_E19_to_W1910_9_0 ;
  wire \net_cnt_lcd_reg[0]_N14_to_S149_9_0 ;
  wire \net_cnt_lcd_reg[0]_S0_G_B3_to_G39_9_0 ;
  wire \net_cnt_lcd_reg[0]_E18_to_W188_7_0 ;
  wire \net_cnt_lcd_reg[0]_S1_G_B4_to_G48_7_0 ;
  wire \net_cnt_lcd_reg[0]_V6S4_to_V6M410_8_0 ;
  wire \net_cnt_lcd_reg[0]_E0_to_W010_9_0 ;
  wire \net_cnt_lcd_reg[0]_S0_F_B3_to_F310_9_0 ;
  wire \net_cnt_lcd_reg[0]_S0_G_B3_to_G310_9_0 ;
  wire \net_cnt_lcd_reg[0]_S22_to_N229_5_0 ;
  wire \net_cnt_lcd_reg[0]_S1_G_B3_to_G39_5_0 ;
  wire \net_cnt_lcd_reg[0]_V6S10_to_V6M1010_5_0 ;
  wire \net_cnt_lcd_reg[0]_S0_G_B3_to_G310_5_0 ;
  wire \net_cnt_lcd_reg[0]_S1_F_B1_to_F17_5_0 ;
  wire \net_cnt_lcd_reg[0]_S0_F_B2_to_F27_5_0 ;
  wire \net_cnt_lcd_reg[0]_S0_G_B1_to_G17_5_0 ;
  wire \net_cnt_lcd_reg[1]_YQ_to_S1_YQ7_5_0 ;
  wire \net_cnt_lcd_reg[1]_V6S4_to_V6M410_5_0 ;
  wire \net_cnt_lcd_reg[1]_H6E5_to_H6M510_8_0 ;
  wire \net_cnt_lcd_reg[1]_S4_to_N411_8_0 ;
  wire \net_cnt_lcd_reg[1]_W9_to_E911_7_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B4_to_G411_7_0 ;
  wire \net_cnt_lcd_reg[1]_S0_to_N08_5_0 ;
  wire \net_cnt_lcd_reg[1]_E20_to_W208_6_0 ;
  wire \net_cnt_lcd_reg[1]_S22_to_N229_6_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B1_to_G19_6_0 ;
  wire \net_cnt_lcd_reg[1]_H6W0_to_LEFT_H6M07_2_0 ;
  wire \net_cnt_lcd_reg[1]_LEFT_V6S2_to_LEFT_V6M210_2_0 ;
  wire \net_cnt_lcd_reg[1]_LEFT_H6A11_to_H6W1110_7_0 ;
  wire \net_cnt_lcd_reg[1]_N20_to_S209_7_0 ;
  wire \net_cnt_lcd_reg[1]_S1_G_B2_to_G29_7_0 ;
  wire \net_cnt_lcd_reg[1]_E2_to_W211_9_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B2_to_G211_9_0 ;
  wire \net_cnt_lcd_reg[1]_V6S8_to_V6M810_5_0 ;
  wire \net_cnt_lcd_reg[1]_E9_to_W910_6_0 ;
  wire \net_cnt_lcd_reg[1]_S1_G_B1_to_G110_6_0 ;
  wire \net_cnt_lcd_reg[1]_H6E0_to_H6M07_8_0 ;
  wire \net_cnt_lcd_reg[1]_S2_to_N28_8_0 ;
  wire \net_cnt_lcd_reg[1]_E22_to_W228_9_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B1_to_G18_9_0 ;
  wire \net_cnt_lcd_reg[1]_E20_to_W207_9_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B2_to_G27_9_0 ;
  wire \net_cnt_lcd_reg[1]_E5_to_W57_6_0 ;
  wire \net_cnt_lcd_reg[1]_S3_to_N38_6_0 ;
  wire \net_cnt_lcd_reg[1]_S3_to_N39_6_0 ;
  wire \net_cnt_lcd_reg[1]_S1_G_B1_to_G19_6_0 ;
  wire \net_cnt_lcd_reg[1]_N5_to_S59_8_0 ;
  wire \net_cnt_lcd_reg[1]_S0_F_B1_to_F19_8_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B3_to_G311_8_0 ;
  wire \net_cnt_lcd_reg[1]_S8_to_N88_5_0 ;
  wire \net_cnt_lcd_reg[1]_S8_to_N89_5_0 ;
  wire \net_cnt_lcd_reg[1]_S1_G_B2_to_G29_5_0 ;
  wire \net_cnt_lcd_reg[1]_W6_to_E610_7_0 ;
  wire \net_cnt_lcd_reg[1]_S1_G_B3_to_G310_7_0 ;
  wire \net_cnt_lcd_reg[1]_E0_to_W010_6_0 ;
  wire \net_cnt_lcd_reg[1]_N23_to_S239_6_0 ;
  wire \net_cnt_lcd_reg[1]_E21_to_W219_7_0 ;
  wire \net_cnt_lcd_reg[1]_S0_F_B1_to_F19_7_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B1_to_G19_7_0 ;
  wire \net_cnt_lcd_reg[1]_E5_to_W57_7_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B1_to_G17_7_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B2_to_G210_5_0 ;
  wire \net_cnt_lcd_reg[1]_S6_to_N68_8_0 ;
  wire \net_cnt_lcd_reg[1]_E11_to_W118_9_0 ;
  wire \net_cnt_lcd_reg[1]_S1_F_B1_to_F18_9_0 ;
  wire \net_cnt_lcd_reg[1]_S1_G_B1_to_G18_9_0 ;
  wire \net_cnt_lcd_reg[1]_S2_to_N211_6_0 ;
  wire \net_cnt_lcd_reg[1]_S0_F_B3_to_F311_6_0 ;
  wire \net_cnt_lcd_reg[1]_S7_to_N711_6_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B2_to_G211_6_0 ;
  wire \net_cnt_lcd_reg[1]_W5_to_E57_10_0 ;
  wire \net_cnt_lcd_reg[1]_S0_F_B1_to_F17_10_0 ;
  wire \net_cnt_lcd_reg[1]_H6E1_to_H6W17_11_0 ;
  wire \net_cnt_lcd_reg[1]_W6_to_E67_10_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B2_to_G27_10_0 ;
  wire \net_cnt_lcd_reg[1]_S6_to_N611_11_0 ;
  wire \net_cnt_lcd_reg[1]_W2_to_E211_10_0 ;
  wire \net_cnt_lcd_reg[1]_S1_F_B4_to_F411_10_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B2_to_G27_5_0 ;
  wire \net_cnt_lcd_reg[1]_E0_to_W011_9_0 ;
  wire \net_cnt_lcd_reg[1]_S1_F_B1_to_F111_9_0 ;
  wire \net_cnt_lcd_reg[1]_S1_G_B1_to_G111_9_0 ;
  wire \net_cnt_lcd_reg[1]_S7_to_N78_10_0 ;
  wire \net_cnt_lcd_reg[1]_S1_F_B1_to_F18_10_0 ;
  wire \net_cnt_lcd_reg[1]_S4_to_N48_11_0 ;
  wire \net_cnt_lcd_reg[1]_W9_to_E98_10_0 ;
  wire \net_cnt_lcd_reg[1]_S1_G_B2_to_G28_10_0 ;
  wire \net_cnt_lcd_reg[1]_S8_to_N88_11_0 ;
  wire \net_cnt_lcd_reg[1]_W13_to_E138_10_0 ;
  wire \net_cnt_lcd_reg[1]_S0_F_B1_to_F18_10_0 ;
  wire \net_cnt_lcd_reg[1]_S0_G_B1_to_G18_10_0 ;
  wire \net_cnt_lcd_reg[1]_V6S0_to_V6M010_8_0 ;
  wire \net_cnt_lcd_reg[1]_E1_to_W110_9_0 ;
  wire \net_cnt_lcd_reg[1]_S1_G_B1_to_G110_9_0 ;
  wire \net_cnt_lcd_reg[1]_S1_F_B1_to_F18_6_0 ;
  wire \net_cnt_lcd_reg[1]_S1_G_B1_to_G18_6_0 ;
  wire \net_cnt_lcd_reg[2]_XQ_to_S0_XQ9_5_0 ;
  wire \net_cnt_lcd_reg[2]_H6E5_to_H6M59_8_0 ;
  wire \net_cnt_lcd_reg[2]_N5_to_S58_8_0 ;
  wire \net_cnt_lcd_reg[2]_S1_F_B2_to_F28_8_0 ;
  wire \net_cnt_lcd_reg[2]_E2_to_W29_6_0 ;
  wire \net_cnt_lcd_reg[2]_S0_to_N010_6_0 ;
  wire \net_cnt_lcd_reg[2]_S0_G_B1_to_G110_6_0 ;
  wire \net_cnt_lcd_reg[2]_V6S4_to_V6M412_8_0 ;
  wire \net_cnt_lcd_reg[2]_N1_to_S111_8_0 ;
  wire \net_cnt_lcd_reg[2]_S1_F_B3_to_F311_8_0 ;
  wire \net_cnt_lcd_reg[2]_S0_G_B3_to_G39_6_0 ;
  wire \net_cnt_lcd_reg[2]_E0_to_W012_9_0 ;
  wire \net_cnt_lcd_reg[2]_N2_to_S211_9_0 ;
  wire \net_cnt_lcd_reg[2]_S0_F_B4_to_F411_9_0 ;
  wire \net_cnt_lcd_reg[2]_E2_to_W29_7_0 ;
  wire \net_cnt_lcd_reg[2]_N1_to_S18_7_0 ;
  wire \net_cnt_lcd_reg[2]_S0_G_B2_to_G28_7_0 ;
  wire \net_cnt_lcd_reg[2]_S1_to_N110_5_0 ;
  wire \net_cnt_lcd_reg[2]_E1_to_W110_6_0 ;
  wire \net_cnt_lcd_reg[2]_S1_G_B3_to_G310_6_0 ;
  wire \net_cnt_lcd_reg[2]_E1_to_W110_7_0 ;
  wire \net_cnt_lcd_reg[2]_S0_F_B4_to_F410_7_0 ;
  wire \net_cnt_lcd_reg[2]_S6_to_N610_11_0 ;
  wire \net_cnt_lcd_reg[2]_W11_to_E1110_10_0 ;
  wire \net_cnt_lcd_reg[2]_S0_F_B3_to_F310_10_0 ;
  wire \net_cnt_lcd_reg[2]_V6N5_to_V6M56_8_0 ;
  wire \net_cnt_lcd_reg[2]_E22_to_W226_9_0 ;
  wire \net_cnt_lcd_reg[2]_S20_to_N207_9_0 ;
  wire \net_cnt_lcd_reg[2]_S0_F_B1_to_F17_9_0 ;
  wire \net_cnt_lcd_reg[2]_S0_G_B1_to_G17_9_0 ;
  wire \net_cnt_lcd_reg[2]_OUT0_to_OUT_W09_6_0 ;
  wire \net_cnt_lcd_reg[2]_S1_G_B3_to_G39_6_0 ;
  wire \net_cnt_lcd_reg[2]_S1_G_B1_to_G110_10_0 ;
  wire \net_cnt_lcd_reg[2]_H6E0_to_H6M09_8_0 ;
  wire \net_cnt_lcd_reg[2]_N4_to_S48_8_0 ;
  wire \net_cnt_lcd_reg[2]_S0_G_B2_to_G28_8_0 ;
  wire \net_cnt_lcd_reg[2]_S1_G_B1_to_G19_5_0 ;
  wire \net_cnt_lcd_reg[2]_S0_G_B2_to_G29_7_0 ;
  wire \net_cnt_lcd_reg[2]_W0_to_E06_7_0 ;
  wire \net_cnt_lcd_reg[2]_S6_to_N67_7_0 ;
  wire \net_cnt_lcd_reg[2]_S0_G_B3_to_G37_7_0 ;
  wire \net_cnt_lcd_reg[2]_S3_to_N310_5_0 ;
  wire \net_cnt_lcd_reg[2]_S0_F_B3_to_F310_5_0 ;
  wire \net_cnt_lcd_reg[2]_S0_G_B4_to_G410_5_0 ;
  wire \net_cnt_lcd_reg[2]_E7_to_W78_9_0 ;
  wire \net_cnt_lcd_reg[2]_S1_F_B4_to_F48_9_0 ;
  wire \net_cnt_lcd_reg[2]_S1_G_B4_to_G48_9_0 ;
  wire \net_cnt_lcd_reg[2]_S1_to_N111_5_0 ;
  wire \net_cnt_lcd_reg[2]_E1_to_W111_6_0 ;
  wire \net_cnt_lcd_reg[2]_S0_F_B4_to_F411_6_0 ;
  wire \net_cnt_lcd_reg[2]_E5_to_W59_9_0 ;
  wire \net_cnt_lcd_reg[2]_E5_to_W59_10_0 ;
  wire \net_cnt_lcd_reg[2]_S0_G_B1_to_G19_10_0 ;
  wire \net_cnt_lcd_reg[2]_V6N0_to_V6M06_5_0 ;
  wire \net_cnt_lcd_reg[2]_H6E0_to_H6W06_11_0 ;
  wire \net_cnt_lcd_reg[2]_W4_to_E46_10_0 ;
  wire \net_cnt_lcd_reg[2]_S10_to_N107_10_0 ;
  wire \net_cnt_lcd_reg[2]_S0_F_B4_to_F47_10_0 ;
  wire \net_cnt_lcd_reg[2]_V6N11_to_V6M116_11_0 ;
  wire \net_cnt_lcd_reg[2]_W18_to_E186_10_0 ;
  wire \net_cnt_lcd_reg[2]_S22_to_N227_10_0 ;
  wire \net_cnt_lcd_reg[2]_S0_G_B1_to_G17_10_0 ;
  wire \net_cnt_lcd_reg[2]_V6S10_to_V6M1012_11_0 ;
  wire \net_cnt_lcd_reg[2]_W1_to_E112_10_0 ;
  wire \net_cnt_lcd_reg[2]_N1_to_S111_10_0 ;
  wire \net_cnt_lcd_reg[2]_S1_F_B1_to_F111_10_0 ;
  wire \net_cnt_lcd_reg[2]_W7_to_E711_9_0 ;
  wire \net_cnt_lcd_reg[2]_S1_F_B2_to_F211_9_0 ;
  wire \net_cnt_lcd_reg[3]_YQ_to_S0_YQ9_5_0 ;
  wire \net_cnt_lcd_reg[3]_V6S2_to_V6M212_5_0 ;
  wire \net_cnt_lcd_reg[3]_H6E2_to_H6M212_8_0 ;
  wire \net_cnt_lcd_reg[3]_N13_to_S1311_8_0 ;
  wire \net_cnt_lcd_reg[3]_S1_F_B4_to_F411_8_0 ;
  wire \net_cnt_lcd_reg[3]_V6S3_to_V6M312_5_0 ;
  wire \net_cnt_lcd_reg[3]_E19_to_W1912_6_0 ;
  wire \net_cnt_lcd_reg[3]_N14_to_S1411_6_0 ;
  wire \net_cnt_lcd_reg[3]_E8_to_W811_7_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B3_to_G311_7_0 ;
  wire \net_cnt_lcd_reg[3]_E14_to_W149_6_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B4_to_G49_6_0 ;
  wire \net_cnt_lcd_reg[3]_V6N5_to_V6M56_5_0 ;
  wire \net_cnt_lcd_reg[3]_H6E5_to_H6M56_8_0 ;
  wire \net_cnt_lcd_reg[3]_S4_to_N47_8_0 ;
  wire \net_cnt_lcd_reg[3]_S1_G_B2_to_G27_8_0 ;
  wire \net_cnt_lcd_reg[3]_H6E7_to_H6M79_8_0 ;
  wire \net_cnt_lcd_reg[3]_N17_to_S178_8_0 ;
  wire \net_cnt_lcd_reg[3]_W23_to_E238_7_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B1_to_G18_7_0 ;
  wire \net_cnt_lcd_reg[3]_S15_to_N1510_5_0 ;
  wire \net_cnt_lcd_reg[3]_E15_to_W1510_6_0 ;
  wire \net_cnt_lcd_reg[3]_S1_G_B2_to_G210_6_0 ;
  wire \net_cnt_lcd_reg[3]_E19_to_W198_9_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B4_to_G48_9_0 ;
  wire \net_cnt_lcd_reg[3]_S18_to_N1810_11_0 ;
  wire \net_cnt_lcd_reg[3]_W16_to_E1610_10_0 ;
  wire \net_cnt_lcd_reg[3]_S0_F_B4_to_F410_10_0 ;
  wire \net_cnt_lcd_reg[3]_V6N2_to_V6M26_5_0 ;
  wire \net_cnt_lcd_reg[3]_H6E2_to_H6M26_8_0 ;
  wire \net_cnt_lcd_reg[3]_S18_to_N187_8_0 ;
  wire \net_cnt_lcd_reg[3]_E14_to_W147_9_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B4_to_G47_9_0 ;
  wire \net_cnt_lcd_reg[3]_OUT1_to_OUT_W19_6_0 ;
  wire \net_cnt_lcd_reg[3]_S1_G_B4_to_G49_6_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B3_to_G38_8_0 ;
  wire \net_cnt_lcd_reg[3]_H6E11_to_H6M119_8_0 ;
  wire \net_cnt_lcd_reg[3]_E23_to_W239_9_0 ;
  wire \net_cnt_lcd_reg[3]_S0_F_B3_to_F39_9_0 ;
  wire \net_cnt_lcd_reg[3]_S16_to_N1610_8_0 ;
  wire \net_cnt_lcd_reg[3]_W21_to_E2110_7_0 ;
  wire \net_cnt_lcd_reg[3]_S1_G_B2_to_G210_7_0 ;
  wire \net_cnt_lcd_reg[3]_H6W6_to_LEFT_H6M69_2_0 ;
  wire \net_cnt_lcd_reg[3]_LEFT_H6B7_to_H6W79_6_0 ;
  wire \net_cnt_lcd_reg[3]_E15_to_W159_7_0 ;
  wire \net_cnt_lcd_reg[3]_S0_F_B3_to_F39_7_0 ;
  wire \net_cnt_lcd_reg[3]_E13_to_W136_6_0 ;
  wire \net_cnt_lcd_reg[3]_E13_to_W136_7_0 ;
  wire \net_cnt_lcd_reg[3]_S11_to_N117_7_0 ;
  wire \net_cnt_lcd_reg[3]_S0_F_B3_to_F37_7_0 ;
  wire \net_cnt_lcd_reg[3]_V6N7_to_V6M76_8_0 ;
  wire \net_cnt_lcd_reg[3]_W12_to_E126_7_0 ;
  wire \net_cnt_lcd_reg[3]_S18_to_N187_7_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B2_to_G27_7_0 ;
  wire \net_cnt_lcd_reg[3]_S17_to_N1710_5_0 ;
  wire \net_cnt_lcd_reg[3]_S0_F_B2_to_F210_5_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B1_to_G110_5_0 ;
  wire \net_cnt_lcd_reg[3]_S1_F_B3_to_F38_9_0 ;
  wire \net_cnt_lcd_reg[3]_S12_to_N1210_6_0 ;
  wire \net_cnt_lcd_reg[3]_S12_to_N1211_6_0 ;
  wire \net_cnt_lcd_reg[3]_S0_F_B2_to_F211_6_0 ;
  wire \net_cnt_lcd_reg[3]_E13_to_W1312_6_0 ;
  wire \net_cnt_lcd_reg[3]_N8_to_S811_6_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B4_to_G411_6_0 ;
  wire \net_cnt_lcd_reg[3]_W23_to_E2310_10_0 ;
  wire \net_cnt_lcd_reg[3]_S21_to_N2111_10_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B2_to_G211_10_0 ;
  wire \net_cnt_lcd_reg[3]_W1_to_E19_10_0 ;
  wire \net_cnt_lcd_reg[3]_S0_F_B3_to_F39_10_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B3_to_G39_10_0 ;
  wire \net_cnt_lcd_reg[3]_V6N7_to_V6M76_11_0 ;
  wire \net_cnt_lcd_reg[3]_W12_to_E126_10_0 ;
  wire \net_cnt_lcd_reg[3]_S18_to_N187_10_0 ;
  wire \net_cnt_lcd_reg[3]_S0_F_B2_to_F27_10_0 ;
  wire \net_cnt_lcd_reg[3]_V6N9_to_V6M96_11_0 ;
  wire \net_cnt_lcd_reg[3]_W6_to_E66_10_0 ;
  wire \net_cnt_lcd_reg[3]_S8_to_N87_10_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B3_to_G37_10_0 ;
  wire \net_cnt_lcd_reg[3]_S1_F_B3_to_F311_10_0 ;
  wire \net_cnt_lcd_reg[3]_N20_to_S208_11_0 ;
  wire \net_cnt_lcd_reg[3]_W22_to_E228_10_0 ;
  wire \net_cnt_lcd_reg[3]_S1_G_B1_to_G18_10_0 ;
  wire \net_cnt_lcd_reg[3]_W15_to_E159_10_0 ;
  wire \net_cnt_lcd_reg[3]_N15_to_S158_10_0 ;
  wire \net_cnt_lcd_reg[3]_S0_F_B3_to_F38_10_0 ;
  wire \net_cnt_lcd_reg[3]_S0_G_B3_to_G38_10_0 ;
  wire \net_cnt_lcd_reg[3]_E12_to_W1210_9_0 ;
  wire \net_cnt_lcd_reg[3]_S1_F_B2_to_F210_9_0 ;
  wire \net_cnt_lcd_reg[3]_S1_G_B2_to_G210_9_0 ;
  wire \net_cnt_lcd_reg[3]_H6W10_to_LEFT_H6M109_2_0 ;
  wire \net_cnt_lcd_reg[3]_LEFT_H6B11_to_H6W119_6_0 ;
  wire \net_cnt_lcd_reg[3]_N20_to_S208_6_0 ;
  wire \net_cnt_lcd_reg[3]_S1_F_B2_to_F28_6_0 ;
  wire \net_cnt_lcd_reg[3]_N18_to_S188_5_0 ;
  wire \net_cnt_lcd_reg[3]_E12_to_W128_6_0 ;
  wire \net_cnt_lcd_reg[3]_S1_G_B3_to_G38_6_0 ;
  wire \net_cnt_lcd_reg[4]_XQ_to_S0_XQ7_6_0 ;
  wire \net_cnt_lcd_reg[4]_S7_to_N78_6_0 ;
  wire \net_cnt_lcd_reg[4]_S7_to_N79_6_0 ;
  wire \net_cnt_lcd_reg[4]_S7_to_N710_6_0 ;
  wire \net_cnt_lcd_reg[4]_S0_F_B4_to_F410_6_0 ;
  wire \net_cnt_lcd_reg[4]_E8_to_W87_7_0 ;
  wire \net_cnt_lcd_reg[4]_E8_to_W87_8_0 ;
  wire \net_cnt_lcd_reg[4]_S0_F_B2_to_F27_8_0 ;
  wire \net_cnt_lcd_reg[4]_H6E1_to_H6W17_12_0 ;
  wire \net_cnt_lcd_reg[4]_V6S1_to_V6M110_12_0 ;
  wire \net_cnt_lcd_reg[4]_H6W1_to_H6M110_9_0 ;
  wire \net_cnt_lcd_reg[4]_S9_to_N911_9_0 ;
  wire \net_cnt_lcd_reg[4]_W10_to_E1011_8_0 ;
  wire \net_cnt_lcd_reg[4]_S1_F_B2_to_F211_8_0 ;
  wire \net_cnt_lcd_reg[4]_V6N1_to_V6M14_6_0 ;
  wire \net_cnt_lcd_reg[4]_V6S2_to_V6N210_6_0 ;
  wire \net_cnt_lcd_reg[4]_S14_to_N1411_6_0 ;
  wire \net_cnt_lcd_reg[4]_E10_to_W1011_7_0 ;
  wire \net_cnt_lcd_reg[4]_S0_G_B2_to_G211_7_0 ;
  wire \net_cnt_lcd_reg[4]_S5_to_N58_6_0 ;
  wire \net_cnt_lcd_reg[4]_S5_to_N59_6_0 ;
  wire \net_cnt_lcd_reg[4]_E5_to_W59_7_0 ;
  wire \net_cnt_lcd_reg[4]_S1_G_B3_to_G39_7_0 ;
  wire \net_cnt_lcd_reg[4]_S1_G_B3_to_G37_8_0 ;
  wire \net_cnt_lcd_reg[4]_S10_to_N108_7_0 ;
  wire \net_cnt_lcd_reg[4]_S0_F_B2_to_F28_7_0 ;
  wire \net_cnt_lcd_reg[4]_S5_to_N510_6_0 ;
  wire \net_cnt_lcd_reg[4]_S1_G_B4_to_G410_6_0 ;
  wire \net_cnt_lcd_reg[4]_S9_to_N98_9_0 ;
  wire \net_cnt_lcd_reg[4]_S0_G_B2_to_G28_9_0 ;
  wire \net_cnt_lcd_reg[4]_H6W1_to_H6M17_3_0 ;
  wire \net_cnt_lcd_reg[4]_V6S1_to_V6M110_3_0 ;
  wire \net_cnt_lcd_reg[4]_H6E1_to_H6W110_9_0 ;
  wire \net_cnt_lcd_reg[4]_W10_to_E1010_8_0 ;
  wire \net_cnt_lcd_reg[4]_S0_F_B3_to_F310_8_0 ;
  wire \net_cnt_lcd_reg[4]_E9_to_W97_10_0 ;
  wire \net_cnt_lcd_reg[4]_S1_F_B1_to_F17_10_0 ;
  wire \net_cnt_lcd_reg[4]_E6_to_W67_10_0 ;
  wire \net_cnt_lcd_reg[4]_S1_G_B2_to_G27_10_0 ;
  wire \net_cnt_lcd_reg[4]_E7_to_W79_7_0 ;
  wire \net_cnt_lcd_reg[4]_S1_to_N110_7_0 ;
  wire \net_cnt_lcd_reg[4]_S0_F_B3_to_F310_7_0 ;
  wire \net_cnt_lcd_reg[4]_E10_to_W1010_7_0 ;
  wire \net_cnt_lcd_reg[4]_S0_G_B2_to_G210_7_0 ;
  wire \net_cnt_lcd_reg[4]_H6E9_to_H6W97_12_0 ;
  wire \net_cnt_lcd_reg[4]_V6S4_to_V6M410_12_0 ;
  wire \net_cnt_lcd_reg[4]_W2_to_E210_11_0 ;
  wire \net_cnt_lcd_reg[4]_W2_to_E210_10_0 ;
  wire \net_cnt_lcd_reg[4]_S0_F_B2_to_F210_10_0 ;
  wire \net_cnt_lcd_reg[4]_S0_G_B1_to_G110_10_0 ;
  wire \net_cnt_lcd_reg[4]_S1_F_B1_to_F19_6_0 ;
  wire \net_cnt_lcd_reg[4]_S1_F_B3_to_F37_7_0 ;
  wire \net_cnt_lcd_reg[4]_W10_to_E108_8_0 ;
  wire \net_cnt_lcd_reg[4]_S12_to_N129_8_0 ;
  wire \net_cnt_lcd_reg[4]_S0_G_B2_to_G29_8_0 ;
  wire \net_cnt_lcd_reg[4]_E7_to_W78_7_0 ;
  wire \net_cnt_lcd_reg[4]_E7_to_W78_8_0 ;
  wire \net_cnt_lcd_reg[4]_S0_F_B2_to_F28_8_0 ;
  wire \net_cnt_lcd_reg[4]_S9_to_N99_9_0 ;
  wire \net_cnt_lcd_reg[4]_S0_F_B2_to_F29_9_0 ;
  wire \net_cnt_lcd_reg[4]_S1_F_B1_to_F18_7_0 ;
  wire \net_cnt_lcd_reg[4]_S1_G_B1_to_G18_7_0 ;
  wire \net_cnt_lcd_reg[4]_S3_to_N310_7_0 ;
  wire \net_cnt_lcd_reg[4]_S1_F_B1_to_F110_7_0 ;
  wire \net_cnt_lcd_reg[4]_S1_G_B1_to_G110_7_0 ;
  wire \net_cnt_lcd_reg[4]_S1_G_B3_to_G38_9_0 ;
  wire \net_cnt_lcd_reg[4]_S0_F_B1_to_F111_6_0 ;
  wire \net_cnt_lcd_reg[4]_S0_G_B1_to_G111_6_0 ;
  wire \net_cnt_lcd_reg[4]_S0_F_B1_to_F18_6_0 ;
  wire \net_cnt_lcd_reg[4]_S1_F_B3_to_F311_7_0 ;
  wire \net_cnt_lcd_reg[4]_S1_G_B3_to_G311_7_0 ;
  wire \net_cnt_lcd_reg[4]_H6W4_to_H6M410_9_0 ;
  wire \net_cnt_lcd_reg[4]_S2_to_N211_9_0 ;
  wire \net_cnt_lcd_reg[4]_E22_to_W2211_10_0 ;
  wire \net_cnt_lcd_reg[4]_S0_G_B1_to_G111_10_0 ;
  wire \net_Lut-U144_0_0_Y_to_S0_Y9_6_0 ;
  wire \net_Lut-U144_0_0_H6E1_to_H6M19_9_0 ;
  wire \net_Lut-U144_0_0_V6N1_to_V6M16_9_0 ;
  wire \net_Lut-U144_0_0_W8_to_E86_8_0 ;
  wire \net_Lut-U144_0_0_S14_to_N147_8_0 ;
  wire \net_Lut-U144_0_0_S0_F_B1_to_F17_8_0 ;
  wire \net_Lut-U144_0_0_E17_to_W179_7_0 ;
  wire \net_Lut-U144_0_0_N12_to_S128_7_0 ;
  wire \net_Lut-U144_0_0_S0_F_B1_to_F18_7_0 ;
  wire \net_Lut-U144_0_0_V6N7_to_V6M76_6_0 ;
  wire \net_Lut-U144_0_0_E10_to_W106_7_0 ;
  wire \net_Lut-U144_0_0_S8_to_N87_7_0 ;
  wire \net_Lut-U144_0_0_S1_F_B2_to_F27_7_0 ;
  wire \net_Lut-U144_0_0_N9_to_S98_6_0 ;
  wire \net_Lut-U144_0_0_S0_F_B2_to_F28_6_0 ;
  wire \net_cnt_lcd_reg[5]_YQ_to_S0_YQ7_6_0 ;
  wire \net_cnt_lcd_reg[5]_V6S4_to_V6M410_6_0 ;
  wire \net_cnt_lcd_reg[5]_E0_to_W010_7_0 ;
  wire \net_cnt_lcd_reg[5]_E0_to_W010_8_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B2_to_F210_8_0 ;
  wire \net_cnt_lcd_reg[5]_H6E5_to_H6M510_9_0 ;
  wire \net_cnt_lcd_reg[5]_N5_to_S59_9_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B4_to_F49_9_0 ;
  wire \net_cnt_lcd_reg[5]_E2_to_W27_7_0 ;
  wire \net_cnt_lcd_reg[5]_E2_to_W27_8_0 ;
  wire \net_cnt_lcd_reg[5]_S0_F_B3_to_F37_8_0 ;
  wire \net_cnt_lcd_reg[5]_S1_to_N18_6_0 ;
  wire \net_cnt_lcd_reg[5]_S1_to_N19_6_0 ;
  wire \net_cnt_lcd_reg[5]_E1_to_W19_7_0 ;
  wire \net_cnt_lcd_reg[5]_S1_G_B1_to_G19_7_0 ;
  wire \net_cnt_lcd_reg[5]_S1_G_B1_to_G17_8_0 ;
  wire \net_cnt_lcd_reg[5]_S4_to_N411_9_0 ;
  wire \net_cnt_lcd_reg[5]_S0_G_B3_to_G311_9_0 ;
  wire \net_cnt_lcd_reg[5]_E1_to_W18_7_0 ;
  wire \net_cnt_lcd_reg[5]_S0_F_B3_to_F38_7_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B2_to_F210_6_0 ;
  wire \net_cnt_lcd_reg[5]_H6E5_to_H6M57_9_0 ;
  wire \net_cnt_lcd_reg[5]_S4_to_N48_9_0 ;
  wire \net_cnt_lcd_reg[5]_S0_G_B3_to_G38_9_0 ;
  wire \net_cnt_lcd_reg[5]_H6E11_to_H6M117_9_0 ;
  wire \net_cnt_lcd_reg[5]_V6S10_to_V6M1010_9_0 ;
  wire \net_cnt_lcd_reg[5]_E21_to_W2110_10_0 ;
  wire \net_cnt_lcd_reg[5]_S0_F_B1_to_F110_10_0 ;
  wire \net_cnt_lcd_reg[5]_H6E0_to_H6M07_9_0 ;
  wire \net_cnt_lcd_reg[5]_S0_G_B3_to_G37_9_0 ;
  wire \net_cnt_lcd_reg[5]_S0_to_N08_6_0 ;
  wire \net_cnt_lcd_reg[5]_S0_to_N09_6_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B4_to_F49_6_0 ;
  wire \net_cnt_lcd_reg[5]_S2_to_N28_6_0 ;
  wire \net_cnt_lcd_reg[5]_S2_to_N29_6_0 ;
  wire \net_cnt_lcd_reg[5]_S1_G_B2_to_G29_6_0 ;
  wire \net_cnt_lcd_reg[5]_E3_to_W37_7_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B1_to_F17_7_0 ;
  wire \net_cnt_lcd_reg[5]_V6S3_to_V6M310_6_0 ;
  wire \net_cnt_lcd_reg[5]_H6E3_to_H6M310_9_0 ;
  wire \net_cnt_lcd_reg[5]_S21_to_N2111_9_0 ;
  wire \net_cnt_lcd_reg[5]_W22_to_E2211_8_0 ;
  wire \net_cnt_lcd_reg[5]_S0_G_B4_to_G411_8_0 ;
  wire \net_cnt_lcd_reg[5]_S17_to_N178_6_0 ;
  wire \net_cnt_lcd_reg[5]_E17_to_W178_7_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B4_to_F48_7_0 ;
  wire \net_cnt_lcd_reg[5]_S0_G_B4_to_G410_9_0 ;
  wire \net_cnt_lcd_reg[5]_E20_to_W209_7_0 ;
  wire \net_cnt_lcd_reg[5]_S0_F_B2_to_F29_7_0 ;
  wire \net_cnt_lcd_reg[5]_OUT0_to_OUT_W07_7_0 ;
  wire \net_cnt_lcd_reg[5]_S0_F_B2_to_F27_7_0 ;
  wire \net_cnt_lcd_reg[5]_W2_to_E210_5_0 ;
  wire \net_cnt_lcd_reg[5]_S0_F_B1_to_F110_5_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B2_to_F28_9_0 ;
  wire \net_cnt_lcd_reg[5]_S1_G_B2_to_G28_9_0 ;
  wire \net_cnt_lcd_reg[5]_V6S0_to_V6M010_6_0 ;
  wire \net_cnt_lcd_reg[5]_S4_to_N411_6_0 ;
  wire \net_cnt_lcd_reg[5]_S0_G_B3_to_G311_6_0 ;
  wire \net_cnt_lcd_reg[5]_V6S4_to_V6M410_9_0 ;
  wire \net_cnt_lcd_reg[5]_E0_to_W010_10_0 ;
  wire \net_cnt_lcd_reg[5]_N23_to_S239_10_0 ;
  wire \net_cnt_lcd_reg[5]_S0_F_B2_to_F29_10_0 ;
  wire \net_cnt_lcd_reg[5]_S0_G_B2_to_G29_10_0 ;
  wire \net_cnt_lcd_reg[5]_E23_to_W237_10_0 ;
  wire \net_cnt_lcd_reg[5]_S0_F_B3_to_F37_10_0 ;
  wire \net_cnt_lcd_reg[5]_E2_to_W27_10_0 ;
  wire \net_cnt_lcd_reg[5]_S0_G_B4_to_G47_10_0 ;
  wire \net_cnt_lcd_reg[5]_H6E0_to_H6M010_9_0 ;
  wire \net_cnt_lcd_reg[5]_S6_to_N611_9_0 ;
  wire \net_cnt_lcd_reg[5]_E2_to_W211_10_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B2_to_F211_10_0 ;
  wire \net_cnt_lcd_reg[5]_S1_G_B2_to_G211_9_0 ;
  wire \net_cnt_lcd_reg[5]_E0_to_W08_10_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B2_to_F28_10_0 ;
  wire \net_cnt_lcd_reg[5]_S6_to_N68_9_0 ;
  wire \net_cnt_lcd_reg[5]_E2_to_W28_10_0 ;
  wire \net_cnt_lcd_reg[5]_S0_F_B2_to_F28_10_0 ;
  wire \net_cnt_lcd_reg[5]_S0_G_B2_to_G28_10_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B1_to_F110_9_0 ;
  wire \net_cnt_lcd_reg[5]_S1_F_B3_to_F38_6_0 ;
  wire \net_cnt_lcd_reg[5]_S1_G_B2_to_G28_6_0 ;
  wire \net_cnt_lcd_reg[7]_YQ_to_S1_YQ7_6_0 ;
  wire \net_cnt_lcd_reg[7]_E15_to_W157_7_0 ;
  wire \net_cnt_lcd_reg[7]_E15_to_W157_8_0 ;
  wire \net_cnt_lcd_reg[7]_E15_to_W157_9_0 ;
  wire \net_cnt_lcd_reg[7]_S1_G_B2_to_G27_9_0 ;
  wire \net_cnt_lcd_reg[7]_E17_to_W177_7_0 ;
  wire \net_cnt_lcd_reg[7]_S15_to_N158_7_0 ;
  wire \net_cnt_lcd_reg[7]_E15_to_W158_8_0 ;
  wire \net_cnt_lcd_reg[7]_S1_G_B2_to_G28_8_0 ;
  wire \net_cnt_lcd_reg[7]_V6S10_to_V6M1010_6_0 ;
  wire \net_cnt_lcd_reg[7]_H6E11_to_H6M1110_9_0 ;
  wire \net_cnt_lcd_reg[7]_S20_to_N2011_9_0 ;
  wire \net_cnt_lcd_reg[7]_S0_F_B1_to_F111_9_0 ;
  wire \net_cnt_lcd_reg[7]_H6E2_to_H6M27_9_0 ;
  wire \net_cnt_lcd_reg[7]_S18_to_N188_9_0 ;
  wire \net_cnt_lcd_reg[7]_S0_F_B2_to_F28_9_0 ;
  wire \net_cnt_lcd_reg[7]_E12_to_W127_10_0 ;
  wire \net_cnt_lcd_reg[7]_S1_F_B2_to_F27_10_0 ;
  wire \net_cnt_lcd_reg[7]_E21_to_W2110_7_0 ;
  wire \net_cnt_lcd_reg[7]_S0_F_B1_to_F110_7_0 ;
  wire \net_cnt_lcd_reg[7]_V6S2_to_V6M210_12_0 ;
  wire \net_cnt_lcd_reg[7]_W15_to_E1510_11_0 ;
  wire \net_cnt_lcd_reg[7]_W15_to_E1510_10_0 ;
  wire \net_cnt_lcd_reg[7]_S0_G_B2_to_G210_10_0 ;
  wire \net_cnt_lcd_reg[7]_S0_F_B2_to_F27_9_0 ;
  wire \net_cnt_lcd_reg[7]_S12_to_N128_6_0 ;
  wire \net_cnt_lcd_reg[7]_S12_to_N129_6_0 ;
  wire \net_cnt_lcd_reg[7]_S1_F_B3_to_F39_6_0 ;
  wire \net_cnt_lcd_reg[7]_V6S6_to_V6M610_6_0 ;
  wire \net_cnt_lcd_reg[7]_H6E7_to_H6M710_9_0 ;
  wire \net_cnt_lcd_reg[7]_E14_to_W1410_10_0 ;
  wire \net_cnt_lcd_reg[7]_S1_F_B1_to_F110_10_0 ;
  wire \net_cnt_lcd_reg[7]_N17_to_S179_9_0 ;
  wire \net_cnt_lcd_reg[7]_S0_G_B1_to_G19_9_0 ;
  wire \net_cnt_lcd_reg[7]_E8_to_W88_7_0 ;
  wire \net_cnt_lcd_reg[7]_S1_F_B2_to_F28_7_0 ;
  wire \net_cnt_lcd_reg[7]_S1_G_B2_to_G28_7_0 ;
  wire \net_cnt_lcd_reg[7]_S0_F_B1_to_F110_9_0 ;
  wire \net_cnt_lcd_reg[7]_S0_G_B1_to_G110_9_0 ;
  wire \net_cnt_lcd_reg[7]_S14_to_N148_6_0 ;
  wire \net_cnt_lcd_reg[7]_S0_G_B1_to_G18_6_0 ;
  wire \net_Lut-U137_0_0_X_to_S0_X8_7_0 ;
  wire \net_Lut-U137_0_0_W21_to_E218_6_0 ;
  wire \net_Lut-U137_0_0_S0_G_B2_to_G28_6_0 ;
  wire \net_Lut-U191_1_Y_to_S0_Y8_7_0 ;
  wire \net_Lut-U191_1_W9_to_E98_6_0 ;
  wire \net_Lut-U191_1_S11_to_N119_6_0 ;
  wire \net_Lut-U191_1_S0_F_B3_to_F39_6_0 ;
  wire \net_Lut-U191_1_N9_to_S97_7_0 ;
  wire \net_Lut-U191_1_S1_G_B1_to_G17_7_0 ;
  wire \net_Lut-U178_0_X_to_S0_X8_8_0 ;
  wire \net_Lut-U178_0_N21_to_S217_8_0 ;
  wire \net_Lut-U178_0_W3_to_E37_7_0 ;
  wire \net_Lut-U178_0_S1_G_B2_to_G27_7_0 ;
  wire \net_Lut-U174_0_X_to_S1_X7_8_0 ;
  wire \net_Lut-U174_0_W11_to_E117_7_0 ;
  wire \net_Lut-U174_0_S1_G_B3_to_G37_7_0 ;
  wire \net_Lut-U126_0_0_Y_to_S1_Y7_8_0 ;
  wire \net_Lut-U126_0_0_S0_G_B1_to_G17_8_0 ;
  wire \net_Lut-U130_0_1_X_to_S1_X7_9_0 ;
  wire \net_Lut-U130_0_1_W23_to_E237_8_0 ;
  wire \net_Lut-U130_0_1_S0_G_B2_to_G27_8_0 ;
  wire \net_Lut-U209_0_0_Y_to_S0_Y8_8_0 ;
  wire \net_Lut-U209_0_0_H6E9_to_H6M98_11_0 ;
  wire \net_Lut-U209_0_0_S8_to_N89_11_0 ;
  wire \net_Lut-U209_0_0_W13_to_E139_10_0 ;
  wire \net_Lut-U209_0_0_S1_G_B3_to_G39_10_0 ;
  wire \net_Lut-U209_0_0_N14_to_S147_8_0 ;
  wire \net_Lut-U209_0_0_S0_G_B3_to_G37_8_0 ;
  wire \net_Lut-U127_0_Y_to_S1_Y7_9_0 ;
  wire \net_Lut-U127_0_OUT6_to_OUT_E67_8_0 ;
  wire \net_Lut-U127_0_S0_G_B4_to_G47_8_0 ;
  wire \net_Lut-U153_0_X_to_S1_X9_9_0 ;
  wire \net_Lut-U153_0_OUT6_to_OUT_E69_8_0 ;
  wire \net_Lut-U153_0_S1_F_B1_to_F19_8_0 ;
  wire \net_Lut-U225_0_X_to_S1_X10_10_0 ;
  wire \net_Lut-U225_0_N9_to_S99_10_0 ;
  wire \net_Lut-U225_0_S1_G_B1_to_G19_10_0 ;
  wire \net_Lut-U225_0_V6N2_to_V6M27_10_0 ;
  wire \net_Lut-U225_0_H6W2_to_H6M27_7_0 ;
  wire \net_Lut-U225_0_S18_to_N188_7_0 ;
  wire \net_Lut-U225_0_E14_to_W148_8_0 ;
  wire \net_Lut-U225_0_S1_F_B1_to_F18_8_0 ;
  wire \net_Lut-U225_0_H6W1_to_H6M110_7_0 ;
  wire \net_Lut-U225_0_W15_to_E1510_6_0 ;
  wire \net_Lut-U225_0_S0_G_B2_to_G210_6_0 ;
  wire \net_Lut-U225_0_H6W2_to_H6M210_7_0 ;
  wire \net_Lut-U225_0_N16_to_S169_7_0 ;
  wire \net_Lut-U225_0_S1_F_B1_to_F19_7_0 ;
  wire \net_Lut-U225_0_N10_to_S109_7_0 ;
  wire \net_Lut-U225_0_E4_to_W49_8_0 ;
  wire \net_Lut-U225_0_S1_F_B2_to_F29_8_0 ;
  wire \net_Lut-U151_0_Y_to_S1_Y9_9_0 ;
  wire \net_Lut-U151_0_W11_to_E119_8_0 ;
  wire \net_Lut-U151_0_S1_F_B3_to_F39_8_0 ;
  wire \net_Lut-U160_0_X_to_S0_X10_8_0 ;
  wire \net_Lut-U160_0_S1_F_B1_to_F110_8_0 ;
  wire \net_Lut-U158_0_Y_to_S0_Y10_8_0 ;
  wire \net_Lut-U158_0_S1_F_B3_to_F310_8_0 ;
  wire \net_Lut-U170_1_X_to_S1_X11_8_0 ;
  wire \net_Lut-U170_1_N12_to_S1210_8_0 ;
  wire \net_Lut-U170_1_S1_F_B4_to_F410_8_0 ;
  wire \net_Lut-U170_1_V6N2_to_V6M28_8_0 ;
  wire \net_Lut-U170_1_S16_to_N169_8_0 ;
  wire \net_Lut-U170_1_S0_F_B2_to_F29_8_0 ;
  wire \net_Lut-U195_0_Y_to_S1_Y10_10_0 ;
  wire \net_Lut-U195_0_W22_to_E2210_9_0 ;
  wire \net_Lut-U195_0_W22_to_E2210_8_0 ;
  wire \net_Lut-U195_0_S1_G_B1_to_G110_8_0 ;
  wire \net_Lut-U196_4_Y_to_S1_Y11_8_0 ;
  wire \net_Lut-U196_4_N0_to_S010_8_0 ;
  wire \net_Lut-U196_4_S1_G_B2_to_G210_8_0 ;
  wire \net_Lut-U196_6_1_X_to_S0_X10_7_0 ;
  wire \net_Lut-U196_6_1_OUT0_to_OUT_W010_8_0 ;
  wire \net_Lut-U196_6_1_S1_G_B3_to_G310_8_0 ;
  wire \net_Lut-U196_7_1_Y_to_S0_Y10_7_0 ;
  wire \net_Lut-U196_7_1_OUT1_to_OUT_W110_8_0 ;
  wire \net_Lut-U196_7_1_S1_G_B4_to_G410_8_0 ;
  wire \net_Lut-U162_0_0_X_to_S0_X9_8_0 ;
  wire \net_Lut-U162_0_0_S1_G_B1_to_G19_8_0 ;
  wire \net_Lut-U165_2_X_to_S1_X9_7_0 ;
  wire \net_Lut-U165_2_E8_to_W89_8_0 ;
  wire \net_Lut-U165_2_S1_G_B2_to_G29_8_0 ;
  wire \net_Lut-U164_0_0_Y_to_S0_Y9_8_0 ;
  wire \net_Lut-U164_0_0_S12_to_N1210_8_0 ;
  wire \net_Lut-U164_0_0_S0_G_B2_to_G210_8_0 ;
  wire \net_Lut-U164_0_0_S1_G_B3_to_G39_8_0 ;
  wire \net_Lut-U115_0_0_Y_to_S1_Y9_7_0 ;
  wire \net_Lut-U115_0_0_W19_to_E199_6_0 ;
  wire \net_Lut-U115_0_0_S0_F_B1_to_F19_6_0 ;
  wire \net_Lut-U121_2_X_to_S0_X10_6_0 ;
  wire \net_Lut-U121_2_N1_to_S19_6_0 ;
  wire \net_Lut-U121_2_S0_F_B2_to_F29_6_0 ;
  wire \net_Lut-U117_0_Y_to_S0_Y10_6_0 ;
  wire \net_Lut-U117_0_N9_to_S99_6_0 ;
  wire \net_Lut-U117_0_S0_F_B4_to_F49_6_0 ;
  wire \net_Lut-U193_0_0_X_to_S1_X8_7_0 ;
  wire \net_Lut-U193_0_0_S0_G_B3_to_G38_7_0 ;
  wire \net_Lut-U213_0_0_Y_to_S1_Y8_7_0 ;
  wire \net_Lut-U213_0_0_S0_G_B4_to_G48_7_0 ;
  wire \net_Lut-U213_0_0_OUT1_to_OUT_W18_8_0 ;
  wire \net_Lut-U213_0_0_S0_G_B1_to_G18_8_0 ;
  wire \net_Lut-U213_0_0_S2_to_N29_7_0 ;
  wire \net_Lut-U213_0_0_S0_G_B3_to_G39_7_0 ;
  wire \net_Lut-U189_2_X_to_S1_X8_8_0 ;
  wire \net_Lut-U189_2_N9_to_S97_8_0 ;
  wire \net_Lut-U189_2_E11_to_W117_9_0 ;
  wire \net_Lut-U189_2_S1_F_B1_to_F17_9_0 ;
  wire \net_Lut-U189_2_S0_F_B1_to_F18_8_0 ;
  wire \net_Lut-U179_2_Y_to_S1_Y8_8_0 ;
  wire \net_Lut-U179_2_S0_F_B3_to_F38_8_0 ;
  wire \net_Lut-U232_0_0_X_to_S0_X7_5_0 ;
  wire \net_Lut-U232_0_0_H6E7_to_H6M77_8_0 ;
  wire \net_Lut-U232_0_0_S16_to_N168_8_0 ;
  wire \net_Lut-U232_0_0_S1_G_B3_to_G38_8_0 ;
  wire \net_Lut-U232_0_0_S1_F_B1_to_F17_8_0 ;
  wire \net_Lut-U232_0_0_V6S6_to_V6M610_5_0 ;
  wire \net_Lut-U232_0_0_H6E7_to_H6M710_8_0 ;
  wire \net_Lut-U232_0_0_S16_to_N1611_8_0 ;
  wire \net_Lut-U232_0_0_E12_to_W1211_9_0 ;
  wire \net_Lut-U232_0_0_S0_F_B2_to_F211_9_0 ;
  wire \net_Lut-U232_0_0_E12_to_W1210_6_0 ;
  wire \net_Lut-U232_0_0_E12_to_W1210_7_0 ;
  wire \net_Lut-U232_0_0_S0_F_B2_to_F210_7_0 ;
  wire \net_Lut-U232_0_0_S15_to_N158_5_0 ;
  wire \net_Lut-U232_0_0_S15_to_N159_5_0 ;
  wire \net_Lut-U232_0_0_E15_to_W159_6_0 ;
  wire \net_Lut-U232_0_0_S1_F_B2_to_F29_6_0 ;
  wire \net_Lut-U232_0_0_S19_to_N198_5_0 ;
  wire \net_Lut-U232_0_0_E19_to_W198_6_0 ;
  wire \net_Lut-U232_0_0_E19_to_W198_7_0 ;
  wire \net_Lut-U232_0_0_S1_F_B3_to_F38_7_0 ;
  wire \net_Lut-U232_0_0_H6W6_to_LEFT_H6M67_2_0 ;
  wire \net_Lut-U232_0_0_LEFT_H6B7_to_H6M77_3_0 ;
  wire \net_Lut-U232_0_0_N17_to_S176_3_0 ;
  wire \net_Lut-U232_0_0_W23_to_LEFT_E236_2_0 ;
  wire \net_Lut-U232_0_0_LEFT_O2_to_OUT6_2_0 ;
  wire \net_Lut-U176_0_1_X_to_S0_X8_9_0 ;
  wire \net_Lut-U176_0_1_N0_to_S07_9_0 ;
  wire \net_Lut-U176_0_1_S1_F_B2_to_F27_9_0 ;
  wire \net_Lut-U176_0_1_S13_to_N139_9_0 ;
  wire \net_Lut-U176_0_1_S1_G_B2_to_G29_9_0 ;
  wire \net_Lut-U176_0_1_N1_to_S17_9_0 ;
  wire \net_Lut-U176_0_1_W7_to_E77_8_0 ;
  wire \net_Lut-U176_0_1_S1_F_B2_to_F27_8_0 ;
  wire \net_Lut-U175_0_0_X_to_S0_X7_7_0 ;
  wire \net_Lut-U175_0_0_OUT0_to_OUT_W07_8_0 ;
  wire \net_Lut-U175_0_0_S1_F_B3_to_F37_8_0 ;
  wire \net_Lut-U204_0_1_Y_to_S0_Y8_9_0 ;
  wire \net_Lut-U204_0_1_S8_to_N89_9_0 ;
  wire \net_Lut-U204_0_1_S1_F_B2_to_F29_9_0 ;
  wire \net_Lut-U204_0_1_W17_to_E178_8_0 ;
  wire \net_Lut-U204_0_1_N17_to_S177_8_0 ;
  wire \net_Lut-U204_0_1_S1_F_B4_to_F47_8_0 ;
  wire \net_Lut-U204_0_1_V6S8_to_V6M811_9_0 ;
  wire \net_Lut-U204_0_1_W13_to_E1311_8_0 ;
  wire \net_Lut-U204_0_1_S0_F_B2_to_F211_8_0 ;
  wire \net_Lut-U204_0_1_S0_G_B2_to_G211_8_0 ;
  wire \net_Lut-U204_0_1_V6S10_to_V6M1011_9_0 ;
  wire \net_Lut-U204_0_1_W1_to_E111_8_0 ;
  wire \net_Lut-U204_0_1_W1_to_E111_7_0 ;
  wire \net_Lut-U204_0_1_S1_F_B2_to_F211_7_0 ;
  wire \net_Lut-U204_0_1_S1_G_B2_to_G211_7_0 ;
  wire \net_Lut-U201_0_0_X_to_S0_X7_9_0 ;
  wire \net_Lut-U201_0_0_W9_to_E97_8_0 ;
  wire \net_Lut-U201_0_0_S11_to_N118_8_0 ;
  wire \net_Lut-U201_0_0_S11_to_N119_8_0 ;
  wire \net_Lut-U201_0_0_W12_to_E129_7_0 ;
  wire \net_Lut-U201_0_0_S1_G_B4_to_G49_7_0 ;
  wire \net_Lut-U201_0_0_W19_to_E197_8_0 ;
  wire \net_Lut-U201_0_0_S1_G_B4_to_G47_8_0 ;
  wire \net_Lut-U201_0_0_V6S0_to_V6M010_9_0 ;
  wire \net_Lut-U201_0_0_W3_to_E310_8_0 ;
  wire \net_Lut-U201_0_0_W3_to_E310_7_0 ;
  wire \net_Lut-U201_0_0_S0_G_B3_to_G310_7_0 ;
  wire \net_Lut-U201_0_0_S0_G_B3_to_G39_8_0 ;
  wire \net_Lut-U201_0_0_V6S1_to_V6M110_9_0 ;
  wire \net_Lut-U201_0_0_W7_to_E710_8_0 ;
  wire \net_Lut-U201_0_0_S5_to_N511_8_0 ;
  wire \net_Lut-U201_0_0_S0_F_B4_to_F411_8_0 ;
  wire \net_Lut-U201_0_0_S1_F_B2_to_F210_7_0 ;
  wire \net_Lut-U201_0_0_W9_to_E97_7_0 ;
  wire \net_Lut-U201_0_0_S0_F_B1_to_F17_7_0 ;
  wire \net_Lut-U201_0_0_V6S8_to_V6M810_9_0 ;
  wire \net_Lut-U201_0_0_W13_to_E1310_8_0 ;
  wire \net_Lut-U201_0_0_W13_to_E1310_7_0 ;
  wire \net_Lut-U201_0_0_S15_to_N1511_7_0 ;
  wire \net_Lut-U201_0_0_S1_F_B4_to_F411_7_0 ;
  wire \net_Lut-U201_0_0_S1_G_B4_to_G411_7_0 ;
  wire \net_Lut-U132_0_Y_to_S0_Y7_9_0 ;
  wire \net_Lut-U132_0_S1_F_B3_to_F37_9_0 ;
  wire \net_Lut-U229_0_X_to_S1_X7_10_0 ;
  wire \net_Lut-U229_0_S5_to_N58_10_0 ;
  wire \net_Lut-U229_0_S5_to_N59_10_0 ;
  wire \net_Lut-U229_0_S1_F_B1_to_F19_10_0 ;
  wire \net_Lut-U229_0_W19_to_E197_9_0 ;
  wire \net_Lut-U229_0_S1_F_B4_to_F47_9_0 ;
  wire \net_Lut-U229_0_S15_to_N158_10_0 ;
  wire \net_Lut-U229_0_W16_to_E168_9_0 ;
  wire \net_Lut-U229_0_S22_to_N229_9_0 ;
  wire \net_Lut-U229_0_S1_G_B4_to_G49_9_0 ;
  wire \net_Lut-U127_0_0_Y_to_S1_Y7_10_0 ;
  wire \net_Lut-U127_0_0_OUT6_to_OUT_E67_9_0 ;
  wire \net_Lut-U127_0_0_S1_G_B1_to_G17_9_0 ;
  wire \net_Lut-U205_0_0_Y_to_S0_Y7_7_0 ;
  wire \net_Lut-U205_0_0_V6S1_to_V6M110_7_0 ;
  wire \net_Lut-U205_0_0_H6E1_to_H6M110_10_0 ;
  wire \net_Lut-U205_0_0_N10_to_S109_10_0 ;
  wire \net_Lut-U205_0_0_W8_to_E89_9_0 ;
  wire \net_Lut-U205_0_0_S1_F_B1_to_F19_9_0 ;
  wire \net_Lut-U205_0_0_S5_to_N58_7_0 ;
  wire \net_Lut-U205_0_0_S5_to_N59_7_0 ;
  wire \net_Lut-U205_0_0_S1_F_B2_to_F29_7_0 ;
  wire \net_Lut-U205_0_0_E7_to_W710_8_0 ;
  wire \net_Lut-U205_0_0_S0_G_B1_to_G110_8_0 ;
  wire \net_Lut-U205_0_0_V6S6_to_V6M610_7_0 ;
  wire \net_Lut-U205_0_0_E12_to_W1210_8_0 ;
  wire \net_Lut-U205_0_0_S14_to_N1411_8_0 ;
  wire \net_Lut-U205_0_0_S0_F_B1_to_F111_8_0 ;
  wire \net_Lut-U205_0_0_S0_G_B1_to_G111_8_0 ;
  wire \net_Lut-U205_0_0_S10_to_N1011_7_0 ;
  wire \net_Lut-U205_0_0_S1_F_B1_to_F111_7_0 ;
  wire \net_Lut-U205_0_0_S5_to_N511_7_0 ;
  wire \net_Lut-U205_0_0_S1_G_B1_to_G111_7_0 ;
  wire \net_Lut-U154_1_X_to_S0_X9_9_0 ;
  wire \net_Lut-U154_1_S1_F_B3_to_F39_9_0 ;
  wire \net_Lut-U227_0_X_to_S1_X10_9_0 ;
  wire \net_Lut-U227_0_E8_to_W810_10_0 ;
  wire \net_Lut-U227_0_N7_to_S79_10_0 ;
  wire \net_Lut-U227_0_S1_F_B3_to_F39_10_0 ;
  wire \net_Lut-U227_0_N9_to_S99_9_0 ;
  wire \net_Lut-U227_0_S1_G_B1_to_G19_9_0 ;
  wire \net_Lut-U152_0_0_X_to_S0_X10_9_0 ;
  wire \net_Lut-U152_0_0_N1_to_S19_9_0 ;
  wire \net_Lut-U152_0_0_S1_G_B3_to_G39_9_0 ;
  wire \net_Lut-U161_0_0_Y_to_S1_Y10_9_0 ;
  wire \net_Lut-U161_0_0_W9_to_E910_8_0 ;
  wire \net_Lut-U161_0_0_S0_F_B1_to_F110_8_0 ;
  wire \net_Lut-U215_0_0_X_to_S1_X11_9_0 ;
  wire \net_Lut-U215_0_0_W7_to_E711_8_0 ;
  wire \net_Lut-U215_0_0_N7_to_S710_8_0 ;
  wire \net_Lut-U215_0_0_S0_F_B2_to_F210_8_0 ;
  wire \net_Lut-U230_0_0_Y_to_S0_Y9_9_0 ;
  wire \net_Lut-U230_0_0_H6W2_to_H6M29_6_0 ;
  wire \net_Lut-U230_0_0_S18_to_N1810_6_0 ;
  wire \net_Lut-U230_0_0_S0_F_B2_to_F210_6_0 ;
  wire \net_Lut-U230_0_0_S15_to_N1510_9_0 ;
  wire \net_Lut-U230_0_0_S15_to_N1511_9_0 ;
  wire \net_Lut-U230_0_0_S0_G_B1_to_G111_9_0 ;
  wire \net_Lut-U230_0_0_W16_to_E1610_8_0 ;
  wire \net_Lut-U230_0_0_S0_F_B4_to_F410_8_0 ;
  wire \net_Lut-U230_0_0_S0_G_B4_to_G410_8_0 ;
  wire \net_Lut-U230_0_0_W17_to_E179_8_0 ;
  wire \net_Lut-U230_0_0_S19_to_N1910_8_0 ;
  wire \net_Lut-U230_0_0_W20_to_E2010_7_0 ;
  wire \net_Lut-U230_0_0_S0_G_B1_to_G110_7_0 ;
  wire \net_Lut-U159_0_0_X_to_S1_X10_7_0 ;
  wire \net_Lut-U159_0_0_E8_to_W810_8_0 ;
  wire \net_Lut-U159_0_0_S0_G_B3_to_G310_8_0 ;
  wire \net_Lut-U170_0_Y_to_S0_Y10_9_0 ;
  wire \net_Lut-U170_0_S12_to_N1211_9_0 ;
  wire \net_Lut-U170_0_W17_to_E1711_8_0 ;
  wire \net_Lut-U170_0_S1_F_B1_to_F111_8_0 ;
  wire \net_Lut-U223_0_X_to_S1_X9_10_0 ;
  wire \net_Lut-U223_0_S8_to_N810_10_0 ;
  wire \net_Lut-U223_0_S1_G_B2_to_G210_10_0 ;
  wire \net_Lut-U208_0_Y_to_S1_Y9_10_0 ;
  wire \net_Lut-U208_0_S17_to_N1710_10_0 ;
  wire \net_Lut-U208_0_S1_G_B3_to_G310_10_0 ;
  wire \net_Lut-U196_1_X_to_S0_X11_7_0 ;
  wire \net_Lut-U196_1_E14_to_W1411_8_0 ;
  wire \net_Lut-U196_1_S1_G_B1_to_G111_8_0 ;
  wire \net_Lut-U196_3_1_Y_to_S0_Y11_7_0 ;
  wire \net_Lut-U196_3_1_E6_to_W611_8_0 ;
  wire \net_Lut-U196_3_1_S1_G_B2_to_G211_8_0 ;
  wire \net_Lut-U196_4_1_X_to_S0_X11_9_0 ;
  wire \net_Lut-U196_4_1_W21_to_E2111_8_0 ;
  wire \net_Lut-U196_4_1_S1_G_B3_to_G311_8_0 ;
  wire \net_Lut-U196_5_1_Y_to_S0_Y11_9_0 ;
  wire \net_Lut-U196_5_1_W9_to_E911_8_0 ;
  wire \net_Lut-U196_5_1_S1_G_B4_to_G411_8_0 ;
  wire \net_Lut-U197_0_0_Y_to_S1_Y10_7_0 ;
  wire \net_Lut-U197_0_0_S13_to_N1311_7_0 ;
  wire \net_Lut-U197_0_0_S0_F_B3_to_F311_7_0 ;
  wire \net_Lut-U197_0_0_S0_G_B4_to_G410_7_0 ;
  wire \net_Lut-U224_0_1_X_to_S0_X9_10_0 ;
  wire \net_Lut-U224_0_1_W9_to_E99_9_0 ;
  wire \net_Lut-U224_0_1_W9_to_E99_8_0 ;
  wire \net_Lut-U224_0_1_S0_F_B3_to_F39_8_0 ;
  wire \net_Lut-U166_0_X_to_S1_X9_6_0 ;
  wire \net_Lut-U166_0_OUT0_to_OUT_W09_7_0 ;
  wire \net_Lut-U166_0_S1_F_B3_to_F39_7_0 ;
  wire \net_Lut-U219_0_1_Y_to_S0_Y9_10_0 ;
  wire \net_Lut-U219_0_1_H6W6_to_H6M69_7_0 ;
  wire \net_Lut-U219_0_1_S1_F_B4_to_F49_7_0 ;
  wire \net_Lut-U190_0_1_X_to_S1_X8_6_0 ;
  wire \net_Lut-U190_0_1_E5_to_W58_7_0 ;
  wire \net_Lut-U190_0_1_E5_to_W58_8_0 ;
  wire \net_Lut-U190_0_1_S1_F_B4_to_F48_8_0 ;
  wire \net_Lut-U190_0_1_E3_to_W38_7_0 ;
  wire \net_Lut-U190_0_1_S21_to_N219_7_0 ;
  wire \net_Lut-U190_0_1_E21_to_W219_8_0 ;
  wire \net_Lut-U190_0_1_S0_G_B1_to_G19_8_0 ;
  wire \net_Lut-U122_0_0_Y_to_S1_Y9_6_0 ;
  wire \net_Lut-U122_0_0_S22_to_N2210_6_0 ;
  wire \net_Lut-U122_0_0_S0_F_B1_to_F110_6_0 ;
  wire \net_Lut-U123_1_X_to_S1_X10_6_0 ;
  wire \net_Lut-U123_1_S0_F_B3_to_F310_6_0 ;
  wire \net_Lut-U186_0_Y_to_S1_Y8_6_0 ;
  wire \net_Lut-U186_0_V6S0_to_V6M011_6_0 ;
  wire \net_Lut-U186_0_N0_to_S010_6_0 ;
  wire \net_Lut-U186_0_S0_G_B3_to_G310_6_0 ;
  wire \net_Lut-U118_0_0_Y_to_S1_Y10_6_0 ;
  wire \net_Lut-U118_0_0_S0_G_B4_to_G410_6_0 ;
  wire \net_Lut-U202_0_0_Y_to_S1_Y11_9_0 ;
  wire \net_Lut-U202_0_0_V6N9_to_V6M98_9_0 ;
  wire \net_Lut-U202_0_0_W6_to_E68_8_0 ;
  wire \net_Lut-U202_0_0_S1_F_B3_to_F38_8_0 ;
  wire \net_Lut-U202_0_0_S0_F_B3_to_F311_9_0 ;
  wire \net_Lut-U202_0_0_OUT7_to_OUT_E711_8_0 ;
  wire \net_Lut-U202_0_0_S0_F_B3_to_F311_8_0 ;
  wire \net_Lut-U180_0_0_X_to_S1_X8_9_0 ;
  wire \net_Lut-U180_0_0_OUT6_to_OUT_E68_8_0 ;
  wire \net_Lut-U180_0_0_S1_G_B1_to_G18_8_0 ;
  wire \net_Lut-U188_0_0_X_to_S0_X8_10_0 ;
  wire \net_Lut-U188_0_0_H6W3_to_H6M38_7_0 ;
  wire \net_Lut-U188_0_0_E21_to_W218_8_0 ;
  wire \net_Lut-U188_0_0_S1_G_B4_to_G48_8_0 ;
  wire \net_Lut-U176_0_0_Y_to_S1_Y8_9_0 ;
  wire \net_Lut-U176_0_0_S0_F_B1_to_F18_9_0 ;
  wire \net_Lut-U177_0_0_X_to_S1_X8_10_0 ;
  wire \net_Lut-U177_0_0_N9_to_S97_10_0 ;
  wire \net_Lut-U177_0_0_S1_G_B1_to_G17_10_0 ;
  wire \net_Lut-U129_0_X_to_S0_X7_10_0 ;
  wire \net_Lut-U129_0_S1_G_B3_to_G37_10_0 ;
  wire \net_Lut-U183_0_0_Y_to_S0_Y8_10_0 ;
  wire \net_Lut-U183_0_0_N12_to_S127_10_0 ;
  wire \net_Lut-U183_0_0_S1_G_B4_to_G47_10_0 ;
  wire \net_Lut-U154_0_Y_to_S0_Y7_10_0 ;
  wire \net_Lut-U154_0_V6S8_to_V6M810_10_0 ;
  wire \net_Lut-U154_0_W13_to_E1310_9_0 ;
  wire \net_Lut-U154_0_N13_to_S139_9_0 ;
  wire \net_Lut-U154_0_S0_F_B1_to_F19_9_0 ;
  wire \net_Lut-U217_1_X_to_S0_X10_10_0 ;
  wire \net_Lut-U217_1_OUT6_to_OUT_E610_9_0 ;
  wire \net_Lut-U217_1_S0_F_B4_to_F410_9_0 ;
  wire \net_Lut-U217_1_S17_to_N1711_10_0 ;
  wire \net_Lut-U217_1_S0_F_B2_to_F211_10_0 ;
  wire \net_Lut-U182_0_1_X_to_S0_X9_7_0 ;
  wire \net_Lut-U182_0_1_S12_to_N1210_7_0 ;
  wire \net_Lut-U182_0_1_S1_F_B3_to_F310_7_0 ;
  wire \net_Lut-U224_0_0_Y_to_S0_Y10_10_0 ;
  wire \net_Lut-U224_0_0_N0_to_S09_10_0 ;
  wire \net_Lut-U224_0_0_S1_F_B2_to_F29_10_0 ;
  wire \net_Lut-U224_0_0_N6_to_S69_10_0 ;
  wire \net_Lut-U224_0_0_S0_F_B1_to_F19_10_0 ;
  wire \net_Lut-U226_0_0_Y_to_S1_Y8_10_0 ;
  wire \net_Lut-U226_0_0_S19_to_N199_10_0 ;
  wire \net_Lut-U226_0_0_S1_F_B4_to_F49_10_0 ;
  wire \net_Lut-U211_0_0_Y_to_S0_Y9_7_0 ;
  wire \net_Lut-U211_0_0_H6E9_to_H6M99_10_0 ;
  wire \net_Lut-U211_0_0_S1_G_B2_to_G29_10_0 ;
  wire \net_Lut-U216_0_X_to_S0_X11_10_0 ;
  wire \net_Lut-U216_0_N13_to_S1310_10_0 ;
  wire \net_Lut-U216_0_N13_to_S139_10_0 ;
  wire \net_Lut-U216_0_S1_G_B4_to_G49_10_0 ;
  wire \net_Lut-U196_0_1_X_to_S0_X11_8_0 ;
  wire \net_Lut-U196_0_1_W16_to_E1611_7_0 ;
  wire \net_Lut-U196_0_1_S0_F_B1_to_F111_7_0 ;
  wire \net_Lut-U196_1_0_Y_to_S0_Y11_8_0 ;
  wire \net_Lut-U196_1_0_W11_to_E1111_7_0 ;
  wire \net_Lut-U196_1_0_S0_F_B2_to_F211_7_0 ;
  wire \net_Lut-U196_2_1_X_to_S1_X11_7_0 ;
  wire \net_Lut-U196_2_1_S0_F_B4_to_F411_7_0 ;
  wire \net_Lut-U196_3_0_Y_to_S1_Y11_7_0 ;
  wire \net_Lut-U196_3_0_S0_G_B1_to_G111_7_0 ;
  wire \net_Lut-U198_0_0_Y_to_S0_Y11_10_0 ;
  wire \net_Lut-U198_0_0_OUT6_to_OUT_E611_9_0 ;
  wire \net_Lut-U198_0_0_S0_G_B4_to_G411_9_0 ;
  wire \net_Lut-U123_0_0_X_to_S0_X10_5_0 ;
  wire \net_Lut-U123_0_0_E11_to_W1110_6_0 ;
  wire \net_Lut-U123_0_0_S1_F_B1_to_F110_6_0 ;
  wire \net_Lut-U124_0_0_X_to_S0_X11_6_0 ;
  wire \net_Lut-U124_0_0_N1_to_S110_6_0 ;
  wire \net_Lut-U124_0_0_S1_F_B3_to_F310_6_0 ;
  wire \net_Lut-U123_2_0_Y_to_S0_Y11_6_0 ;
  wire \net_Lut-U123_2_0_N13_to_S1310_6_0 ;
  wire \net_Lut-U123_2_0_S1_F_B4_to_F410_6_0 ;
  wire \net_Lut-U216_0_0_X_to_S1_X11_10_0 ;
  wire \net_Lut-U216_0_0_S0_F_B1_to_F111_10_0 ;
  wire net_U113_Y_to_S1_Y11_10_0;
  wire net_U113_H6W8_to_H6E811_4_0;
  wire net_U113_V6N9_to_V6M98_4_0;
  wire net_U113_W6_to_E68_3_0;
  wire net_U113_N10_to_S107_3_0;
  wire net_U113_S0_F_B2_to_F27_3_0;
  wire net_U113_S0_G_B2_to_G27_3_0;
  wire net_U113_H6W1_to_H6E111_4_0;
  wire net_U113_W6_to_E611_3_0;
  wire net_U113_N10_to_S1010_3_0;
  wire net_U113_N10_to_S109_3_0;
  wire net_U113_S0_F_B2_to_F29_3_0;
  wire net_U113_S0_G_B2_to_G29_3_0;
  wire net_U113_V6N2_to_V6M28_4_0;
  wire net_U113_S16_to_N169_4_0;
  wire net_U113_S0_F_B2_to_F29_4_0;
  wire net_U113_S0_G_B2_to_G29_4_0;
  wire net_U113_H6W2_to_H6M211_7_0;
  wire net_U113_V6N2_to_V6M28_7_0;
  wire net_U113_W15_to_E158_6_0;
  wire net_U113_N15_to_S157_6_0;
  wire net_U113_S1_F_B2_to_F27_6_0;
  wire net_U113_S1_G_B2_to_G27_6_0;
  wire net_U113_N6_to_S610_4_0;
  wire net_U113_E0_to_W010_5_0;
  wire net_U113_N23_to_S239_5_0;
  wire net_U113_S0_F_B2_to_F29_5_0;
  wire net_U113_S0_G_B2_to_G29_5_0;
  wire net_U113_H6W4_to_H6M411_7_0;
  wire net_U113_V6N5_to_V6M58_7_0;
  wire net_U113_W0_to_E08_6_0;
  wire net_U113_N4_to_S47_6_0;
  wire net_U113_S0_F_B2_to_F27_6_0;
  wire net_U113_S0_G_B2_to_G27_6_0;
  wire net_U113_E13_to_W138_5_0;
  wire net_U113_S11_to_N119_5_0;
  wire net_U113_S1_F_B2_to_F29_5_0;
  wire net_U113_V6N3_to_V6M38_4_0;
  wire net_U113_E19_to_W198_5_0;
  wire net_U113_N14_to_S147_5_0;
  wire net_U113_S1_F_B2_to_F27_5_0;
  wire net_U113_S1_G_B2_to_G27_5_0;
  wire net_U113_W15_to_E158_3_0;
  wire net_U113_S13_to_N139_3_0;
  wire net_U113_S1_F_B2_to_F29_3_0;
  wire net_U113_W21_to_E215_3_0;
  wire net_U113_S23_to_N236_3_0;
  wire net_U113_W0_to_LEFT_E06_2_0;
  wire net_U113_LEFT_O1_to_OUT6_2_0;
  wire \net_Buf-pad-rst_n_IN_to_RIGHT_I35_54_0 ;
  wire \net_Buf-pad-rst_n_RIGHT_LLH2_to_LLH05_5_0 ;
  wire \net_Buf-pad-rst_n_V6S1_to_V6M18_5_0 ;
  wire \net_Buf-pad-rst_n_S5_to_N59_5_0 ;
  wire \net_Buf-pad-rst_n_S1_F_B1_to_F19_5_0 ;
  wire \net_Buf-pad-rst_n_RIGHT_LLH3_to_LLH05_6_0 ;
  wire \net_Buf-pad-rst_n_H6W1_to_H6M15_3_0 ;
  wire \net_Buf-pad-rst_n_V6S1_to_V6N111_3_0 ;
  wire \net_Buf-pad-rst_n_S10_to_N1012_3_0 ;
  wire \net_Buf-pad-rst_n_S10_to_N1013_3_0 ;
  wire \net_Buf-pad-rst_n_W15_to_LEFT_E1513_2_0 ;
  wire \net_Buf-pad-rst_n_LEFT_O3_to_OUT13_2_0 ;
  wire \net_Lut-U149_0_Y_to_S0_Y7_5_0 ;
  wire \net_Lut-U149_0_S1_G_B1_to_G17_5_0 ;
  wire \net_Lut-U147_0_Y_to_S1_Y9_5_0 ;
  wire \net_Lut-U147_0_S0_F_B1_to_F19_5_0 ;
  wire \net_Lut-U145_0_Y_to_S0_Y10_5_0 ;
  wire \net_Lut-U145_0_N13_to_S139_5_0 ;
  wire \net_Lut-U145_0_S0_G_B1_to_G19_5_0 ;
  wire \net_Lut-U143_0_X_to_S0_X8_6_0 ;
  wire \net_Lut-U143_0_N6_to_S67_6_0 ;
  wire \net_Lut-U143_0_S0_F_B1_to_F17_6_0 ;
  wire \net_Lut-U141_0_X_to_S1_X7_7_0 ;
  wire \net_Lut-U141_0_W10_to_E107_6_0 ;
  wire \net_Lut-U141_0_S0_G_B1_to_G17_6_0 ;
  wire \net_Lut-U138_0_X_to_S0_X7_8_0 ;
  wire \net_Lut-U138_0_W19_to_E197_7_0 ;
  wire \net_Lut-U138_0_W19_to_E197_6_0 ;
  wire \net_Lut-U138_0_S1_F_B1_to_F17_6_0 ;
  wire \net_Lut-U136_0_Y_to_S0_Y8_6_0 ;
  wire \net_Lut-U136_0_N9_to_S97_6_0 ;
  wire \net_Lut-U136_0_S1_G_B1_to_G17_6_0 ;
  wire \net_Lut-U173_1_Y_to_S1_Y7_7_0 ;
  wire \net_Lut-U173_1_H6W6_to_H6M67_4_0 ;
  wire \net_Lut-U173_1_W12_to_E127_3_0 ;
  wire \net_Lut-U173_1_S0_F_B1_to_F17_3_0 ;
  wire \net_Lut-U126_1_Y_to_S0_Y7_8_0 ;
  wire \net_Lut-U126_1_H6W10_to_LEFT_H6E107_2_0 ;
  wire \net_Lut-U126_1_LEFT_H6D11_to_H6W117_3_0 ;
  wire \net_Lut-U126_1_S0_G_B1_to_G17_3_0 ;
  wire \net_Lut-U150_0_X_to_S1_X9_8_0 ;
  wire \net_Lut-U150_0_H6W10_to_LEFT_H6E109_2_0 ;
  wire \net_Lut-U150_0_LEFT_H6D11_to_H6W119_3_0 ;
  wire \net_Lut-U150_0_S0_F_B1_to_F19_3_0 ;
  wire \net_Lut-U157_1_X_to_S1_X10_8_0 ;
  wire \net_Lut-U157_1_H6W10_to_LEFT_H6E1010_2_0 ;
  wire \net_Lut-U157_1_LEFT_H6D11_to_H6W1110_3_0 ;
  wire \net_Lut-U157_1_N20_to_S209_3_0 ;
  wire \net_Lut-U157_1_S0_G_B1_to_G19_3_0 ;
  wire \net_Lut-U195_1_Y_to_S1_Y10_8_0 ;
  wire \net_Lut-U195_1_H6W3_to_H6M310_5_0 ;
  wire \net_Lut-U195_1_N22_to_S229_5_0 ;
  wire \net_Lut-U195_1_W20_to_E209_4_0 ;
  wire \net_Lut-U195_1_S0_F_B1_to_F19_4_0 ;
  wire \net_Lut-U162_1_Y_to_S1_Y9_8_0 ;
  wire \net_Lut-U162_1_H6W6_to_H6M69_5_0 ;
  wire \net_Lut-U162_1_W12_to_E129_4_0 ;
  wire \net_Lut-U162_1_S0_G_B1_to_G19_4_0 ;
  wire \net_Lut-U115_1_X_to_S0_X9_6_0 ;
  wire \net_Lut-U115_1_H6W8_to_H6M89_3_0 ;
  wire \net_Lut-U115_1_S1_F_B1_to_F19_3_0 ;
  wire \net_Buf-pad-clk_GCLKOUT_to_CLKB_CLKPAD135_28_0 ;
  wire \net_Buf-pad-clk_CLKB_GCLKBUF1_IN_to_IN35_28_0 ;
  wire net_U108_X_to_S0_X6_3_0;
  wire net_U108_V6S8_to_V6N812_3_0;
  wire net_U108_S5_to_N513_3_0;
  wire net_U108_S5_to_N514_3_0;
  wire net_U108_W6_to_LEFT_E614_2_0;
  wire net_U108_LEFT_O1_to_OUT14_2_0;
  wire net_U108_N12_to_S125_3_0;
  wire net_U108_W14_to_LEFT_E145_2_0;
  wire net_U108_LEFT_O3_to_OUT5_2_0;
  wire \net_lcd_db_reg[6]_XQ_to_S0_XQ9_3_0 ;
  wire \net_lcd_db_reg[6]_OUT7_to_LEFT_OUT_E79_2_0 ;
  wire \net_lcd_db_reg[6]_LEFT_O2_to_OUT9_2_0 ;
  wire \net_lcd_db_reg[5]_YQ_to_S0_YQ9_3_0 ;
  wire \net_lcd_db_reg[5]_W16_to_LEFT_E169_2_0 ;
  wire \net_lcd_db_reg[5]_LEFT_O3_to_OUT9_2_0 ;
  wire \net_lcd_db_reg[4]_YQ_to_S0_YQ9_4_0 ;
  wire \net_lcd_db_reg[4]_W11_to_E119_3_0 ;
  wire \net_lcd_db_reg[4]_S9_to_N910_3_0 ;
  wire \net_lcd_db_reg[4]_W10_to_LEFT_E1010_2_0 ;
  wire \net_lcd_db_reg[4]_LEFT_O1_to_OUT10_2_0 ;
  wire \net_lcd_db_reg[3]_XQ_to_S0_XQ7_3_0 ;
  wire \net_lcd_db_reg[3]_V6S2_to_V6M210_3_0 ;
  wire \net_lcd_db_reg[3]_W15_to_LEFT_E1510_2_0 ;
  wire \net_lcd_db_reg[3]_LEFT_O2_to_OUT10_2_0 ;
  wire \net_lcd_db_reg[2]_XQ_to_S0_XQ9_4_0 ;
  wire \net_lcd_db_reg[2]_N8_to_S88_4_0 ;
  wire \net_lcd_db_reg[2]_W10_to_E108_3_0 ;
  wire \net_lcd_db_reg[2]_W10_to_LEFT_E108_2_0 ;
  wire \net_lcd_db_reg[2]_LEFT_O1_to_OUT8_2_0 ;
  wire \net_lcd_db_reg[1]_XQ_to_S1_XQ9_3_0 ;
  wire \net_lcd_db_reg[1]_W11_to_LEFT_E119_2_0 ;
  wire \net_lcd_db_reg[1]_LEFT_O1_to_OUT9_2_0 ;
  wire \net_lcd_db_reg[0]_YQ_to_S0_YQ7_3_0 ;
  wire \net_lcd_db_reg[0]_V6N1_to_V6M14_3_0 ;
  wire \net_lcd_db_reg[0]_W8_to_LEFT_E84_2_0 ;
  wire \net_lcd_db_reg[0]_LEFT_O1_to_OUT4_2_0 ;
  wire \net_IBuf-clkpad-clk_OUT_to_CLKB_GCLK1_PW35_28_0 ;
  wire \net_IBuf-clkpad-clk_CLKB_GCLK1_to_CLKC_GCLK118_28_0 ;
  wire \net_IBuf-clkpad-clk_CLKC_HGCLK1_to_BRAM_CLKH_GCLK118_1_0 ;
  wire \net_IBuf-clkpad-clk_BRAM_CLKH_VGCLK1_to_BRAM_GCLKIN17_1_0 ;
  wire \net_IBuf-clkpad-clk_BRAM_GCLK_CLBB1_to_GCLK17_3_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK7_3_0 ;
  wire \net_IBuf-clkpad-clk_BRAM_GCLK_CLBD1_to_GCLK19_3_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK9_3_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK9_4_0 ;
  wire \net_IBuf-clkpad-clk_S1_CLK_B_to_CLK7_6_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK9_5_0 ;
  wire \net_IBuf-clkpad-clk_S0_CLK_B_to_CLK7_6_0 ;
  wire \net_IBuf-clkpad-clk_S1_CLK_B_to_CLK7_5_0 ;
  wire \net_IBuf-clkpad-clk_S1_CLK_B_to_CLK9_3_0 ;
  wire net_rst_nInvLut_X_to_S1_X9_5_0;
  wire net_rst_nInvLut_V6N9_to_V6M96_5_0;
  wire net_rst_nInvLut_H6W8_to_LEFT_H6M86_2_0;
  wire net_rst_nInvLut_LEFT_H6B9_to_H6M96_3_0;
  wire net_rst_nInvLut_S8_to_N87_3_0;
  wire net_rst_nInvLut_S0_SR_B_to_SR7_3_0;
  wire net_rst_nInvLut_W10_to_E109_4_0;
  wire net_rst_nInvLut_W10_to_E109_3_0;
  wire net_rst_nInvLut_S0_SR_B_to_SR9_3_0;
  wire net_rst_nInvLut_S0_SR_B_to_SR9_4_0;
  wire net_rst_nInvLut_V6N7_to_V6M76_5_0;
  wire net_rst_nInvLut_E10_to_W106_6_0;
  wire net_rst_nInvLut_S8_to_N87_6_0;
  wire net_rst_nInvLut_S1_SR_B_to_SR7_6_0;
  wire net_rst_nInvLut_S0_SR_B_to_SR9_5_0;
  wire net_rst_nInvLut_S0_SR_B_to_SR7_6_0;
  wire net_rst_nInvLut_V6N1_to_V6B17_5_0;
  wire net_rst_nInvLut_S1_SR_B_to_SR7_5_0;
  wire net_rst_nInvLut_S1_SR_B_to_SR9_3_0;


  defparam iSlice__0___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*~A2)*A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*A1)";
  defparam iSlice__0___inst.fxmux.CONF = "F";
  defparam iSlice__0___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*A1)";
  defparam iSlice__0___inst.gymux.CONF = "G";
  defparam iSlice__0___inst.xused.CONF = "0";
  defparam iSlice__0___inst.yused.CONF = "0";
  defparam iSlice__0___inst.f.INIT = 16'heae0;
  defparam iSlice__0___inst.g.INIT = 16'hfcfe;
  SLICE iSlice__0___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U229_0_S1_F_B1_to_F19_10_0 ),
    .F2(\net_Lut-U224_0_0_S1_F_B2_to_F29_10_0 ),
    .F3(\net_Lut-U227_0_S1_F_B3_to_F39_10_0 ),
    .F4(\net_Lut-U226_0_0_S1_F_B4_to_F49_10_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U225_0_S1_G_B1_to_G19_10_0 ),
    .G2(\net_Lut-U211_0_0_S1_G_B2_to_G29_10_0 ),
    .G3(\net_Lut-U209_0_0_S1_G_B3_to_G39_10_0 ),
    .G4(\net_Lut-U216_0_S1_G_B4_to_G49_10_0 ),
    .XQ(),
    .X(\net_Lut-U223_0_X_to_S1_X9_10_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U208_0_Y_to_S1_Y9_10_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__1___inst.f.CONF = "#LUT:D=(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__1___inst.fxmux.CONF = "F";
  defparam iSlice__1___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*~A2)*A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*~A2)*A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*~A2)*A1)+(((~A4*~A3)*~A2)*A1)";
  defparam iSlice__1___inst.gymux.CONF = "G";
  defparam iSlice__1___inst.xused.CONF = "0";
  defparam iSlice__1___inst.yused.CONF = "0";
  defparam iSlice__1___inst.f.INIT = 16'h7;
  defparam iSlice__1___inst.g.INIT = 16'haaa2;
  SLICE iSlice__1___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U160_0_S1_F_B1_to_F110_8_0 ),
    .F2(\net_cnt_lcd_reg[5]_S1_F_B2_to_F210_8_0 ),
    .F3(\net_Lut-U158_0_S1_F_B3_to_F310_8_0 ),
    .F4(\net_Lut-U170_1_S1_F_B4_to_F410_8_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U195_0_S1_G_B1_to_G110_8_0 ),
    .G2(\net_Lut-U196_4_S1_G_B2_to_G210_8_0 ),
    .G3(\net_Lut-U196_6_1_S1_G_B3_to_G310_8_0 ),
    .G4(\net_Lut-U196_7_1_S1_G_B4_to_G410_8_0 ),
    .XQ(),
    .X(\net_Lut-U157_1_X_to_S1_X10_8_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U195_1_Y_to_S1_Y10_8_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__2___inst.f.CONF = "#LUT:D=(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__2___inst.fxmux.CONF = "F";
  defparam iSlice__2___inst.g.CONF = "#LUT:D=(((A4*~A3)*~A2)*~A1)";
  defparam iSlice__2___inst.gymux.CONF = "G";
  defparam iSlice__2___inst.xused.CONF = "0";
  defparam iSlice__2___inst.yused.CONF = "0";
  defparam iSlice__2___inst.f.INIT = 16'h111;
  defparam iSlice__2___inst.g.INIT = 16'h100;
  SLICE iSlice__2___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U189_2_S1_F_B1_to_F17_9_0 ),
    .F2(\net_Lut-U176_0_1_S1_F_B2_to_F27_9_0 ),
    .F3(\net_Lut-U132_0_S1_F_B3_to_F37_9_0 ),
    .F4(\net_Lut-U229_0_S1_F_B4_to_F47_9_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U127_0_0_S1_G_B1_to_G17_9_0 ),
    .G2(\net_cnt_lcd_reg[7]_S1_G_B2_to_G27_9_0 ),
    .G3(\net_cnt_lcd_reg[6]_S1_G_B3_to_G37_9_0 ),
    .G4(\net_cnt_lcd_reg[0]_S1_G_B4_to_G47_9_0 ),
    .XQ(),
    .X(\net_Lut-U130_0_1_X_to_S1_X7_9_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U127_0_Y_to_S1_Y7_9_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__3___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*A2)*~A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__3___inst.fxmux.CONF = "F";
  defparam iSlice__3___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)";
  defparam iSlice__3___inst.gymux.CONF = "G";
  defparam iSlice__3___inst.xused.CONF = "0";
  defparam iSlice__3___inst.yused.CONF = "0";
  defparam iSlice__3___inst.f.INIT = 16'hefcf;
  defparam iSlice__3___inst.g.INIT = 16'hfefc;
  SLICE iSlice__3___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U205_0_0_S1_F_B1_to_F19_9_0 ),
    .F2(\net_Lut-U204_0_1_S1_F_B2_to_F29_9_0 ),
    .F3(\net_Lut-U154_1_S1_F_B3_to_F39_9_0 ),
    .F4(\net_cnt_lcd_reg[5]_S1_F_B4_to_F49_9_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U227_0_S1_G_B1_to_G19_9_0 ),
    .G2(\net_Lut-U176_0_1_S1_G_B2_to_G29_9_0 ),
    .G3(\net_Lut-U152_0_0_S1_G_B3_to_G39_9_0 ),
    .G4(\net_Lut-U229_0_S1_G_B4_to_G49_9_0 ),
    .XQ(),
    .X(\net_Lut-U153_0_X_to_S1_X9_9_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U151_0_Y_to_S1_Y9_9_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__4___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*~A2)*A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*~A2)*A1)+(((~A4*A3)*A2)*A1)";
  defparam iSlice__4___inst.fxmux.CONF = "F";
  defparam iSlice__4___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*~A1)+(((~A4*A3)*~A2)*~A1)";
  defparam iSlice__4___inst.gymux.CONF = "G";
  defparam iSlice__4___inst.xused.CONF = "0";
  defparam iSlice__4___inst.yused.CONF = "0";
  defparam iSlice__4___inst.f.INIT = 16'haa80;
  defparam iSlice__4___inst.g.INIT = 16'hd010;
  SLICE iSlice__4___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U225_0_S1_F_B1_to_F18_8_0 ),
    .F2(\net_cnt_lcd_reg[2]_S1_F_B2_to_F28_8_0 ),
    .F3(\net_Lut-U202_0_0_S1_F_B3_to_F38_8_0 ),
    .F4(\net_Lut-U190_0_1_S1_F_B4_to_F48_8_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U180_0_0_S1_G_B1_to_G18_8_0 ),
    .G2(\net_cnt_lcd_reg[7]_S1_G_B2_to_G28_8_0 ),
    .G3(\net_Lut-U232_0_0_S1_G_B3_to_G38_8_0 ),
    .G4(\net_Lut-U188_0_0_S1_G_B4_to_G48_8_0 ),
    .XQ(),
    .X(\net_Lut-U189_2_X_to_S1_X8_8_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U179_2_Y_to_S1_Y8_8_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__5___inst.f.CONF = "#LUT:D=(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((~A4*A3)*A2)*~A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)";
  defparam iSlice__5___inst.fxmux.CONF = "F";
  defparam iSlice__5___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*~A2)*A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__5___inst.gymux.CONF = "G";
  defparam iSlice__5___inst.xused.CONF = "0";
  defparam iSlice__5___inst.yused.CONF = "0";
  defparam iSlice__5___inst.f.INIT = 16'hc4c;
  defparam iSlice__5___inst.g.INIT = 16'h7f33;
  SLICE iSlice__5___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U122_0_0_S0_F_B1_to_F110_6_0 ),
    .F2(\net_Lut-U230_0_0_S0_F_B2_to_F210_6_0 ),
    .F3(\net_Lut-U123_1_S0_F_B3_to_F310_6_0 ),
    .F4(\net_cnt_lcd_reg[4]_S0_F_B4_to_F410_6_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[2]_S0_G_B1_to_G110_6_0 ),
    .G2(\net_Lut-U225_0_S0_G_B2_to_G210_6_0 ),
    .G3(\net_Lut-U186_0_S0_G_B3_to_G310_6_0 ),
    .G4(\net_Lut-U118_0_0_S0_G_B4_to_G410_6_0 ),
    .XQ(),
    .X(\net_Lut-U121_2_X_to_S0_X10_6_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U117_0_Y_to_S0_Y10_6_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__6___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__6___inst.fxmux.CONF = "F";
  defparam iSlice__6___inst.g.CONF = "#LUT:D=(((~A4*~A3)*A2)*~A1)";
  defparam iSlice__6___inst.gymux.CONF = "G";
  defparam iSlice__6___inst.xused.CONF = "0";
  defparam iSlice__6___inst.yused.CONF = "0";
  defparam iSlice__6___inst.f.INIT = 16'h807f;
  defparam iSlice__6___inst.g.INIT = 16'h4;
  SLICE iSlice__6___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U144_0_0_S0_F_B1_to_F17_8_0 ),
    .F2(\net_cnt_lcd_reg[4]_S0_F_B2_to_F27_8_0 ),
    .F3(\net_cnt_lcd_reg[5]_S0_F_B3_to_F37_8_0 ),
    .F4(\net_cnt_lcd_reg[6]_S0_F_B4_to_F47_8_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U126_0_0_S0_G_B1_to_G17_8_0 ),
    .G2(\net_Lut-U130_0_1_S0_G_B2_to_G27_8_0 ),
    .G3(\net_Lut-U209_0_0_S0_G_B3_to_G37_8_0 ),
    .G4(\net_Lut-U127_0_S0_G_B4_to_G47_8_0 ),
    .XQ(),
    .X(\net_Lut-U138_0_X_to_S0_X7_8_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U126_1_Y_to_S0_Y7_8_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__7___inst.f.CONF = "#LUT:D=(((A4*~A3)*~A2)*A1)+(((~A4*A3)*A2)*A1)+(((~A4*~A3)*A2)*A1)";
  defparam iSlice__7___inst.fxmux.CONF = "F";
  defparam iSlice__7___inst.g.CONF = "#LUT:D=(((~A4*~A3)*~A2)*A1)";
  defparam iSlice__7___inst.gymux.CONF = "G";
  defparam iSlice__7___inst.xused.CONF = "0";
  defparam iSlice__7___inst.yused.CONF = "0";
  defparam iSlice__7___inst.f.INIT = 16'h288;
  defparam iSlice__7___inst.g.INIT = 16'h2;
  SLICE iSlice__7___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U170_0_S1_F_B1_to_F111_8_0 ),
    .F2(\net_cnt_lcd_reg[4]_S1_F_B2_to_F211_8_0 ),
    .F3(\net_cnt_lcd_reg[2]_S1_F_B3_to_F311_8_0 ),
    .F4(\net_cnt_lcd_reg[3]_S1_F_B4_to_F411_8_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U196_1_S1_G_B1_to_G111_8_0 ),
    .G2(\net_Lut-U196_3_1_S1_G_B2_to_G211_8_0 ),
    .G3(\net_Lut-U196_4_1_S1_G_B3_to_G311_8_0 ),
    .G4(\net_Lut-U196_5_1_S1_G_B4_to_G411_8_0 ),
    .XQ(),
    .X(\net_Lut-U170_1_X_to_S1_X11_8_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U196_4_Y_to_S1_Y11_8_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__8___inst.f.CONF = "#LUT:D=(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__8___inst.fxmux.CONF = "F";
  defparam iSlice__8___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*~A2)*A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*~A2)*A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*~A2)*A1)+(((~A4*~A3)*~A2)*A1)";
  defparam iSlice__8___inst.gymux.CONF = "G";
  defparam iSlice__8___inst.xused.CONF = "0";
  defparam iSlice__8___inst.yused.CONF = "0";
  defparam iSlice__8___inst.f.INIT = 16'h51;
  defparam iSlice__8___inst.g.INIT = 16'haaa2;
  SLICE iSlice__8___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U196_0_1_S0_F_B1_to_F111_7_0 ),
    .F2(\net_Lut-U196_1_0_S0_F_B2_to_F211_7_0 ),
    .F3(\net_Lut-U197_0_0_S0_F_B3_to_F311_7_0 ),
    .F4(\net_Lut-U196_2_1_S0_F_B4_to_F411_7_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U196_3_0_S0_G_B1_to_G111_7_0 ),
    .G2(\net_cnt_lcd_reg[4]_S0_G_B2_to_G211_7_0 ),
    .G3(\net_cnt_lcd_reg[3]_S0_G_B3_to_G311_7_0 ),
    .G4(\net_cnt_lcd_reg[1]_S0_G_B4_to_G411_7_0 ),
    .XQ(),
    .X(\net_Lut-U196_1_X_to_S0_X11_7_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U196_3_1_Y_to_S0_Y11_7_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__9___inst.f.CONF = "#LUT:D=(((A4*~A3)*~A2)*~A1)";
  defparam iSlice__9___inst.fxmux.CONF = "F";
  defparam iSlice__9___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)";
  defparam iSlice__9___inst.gymux.CONF = "G";
  defparam iSlice__9___inst.xused.CONF = "0";
  defparam iSlice__9___inst.yused.CONF = "0";
  defparam iSlice__9___inst.f.INIT = 16'h100;
  defparam iSlice__9___inst.g.INIT = 16'h8000;
  SLICE iSlice__9___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U115_0_0_S0_F_B1_to_F19_6_0 ),
    .F2(\net_Lut-U121_2_S0_F_B2_to_F29_6_0 ),
    .F3(\net_Lut-U191_1_S0_F_B3_to_F39_6_0 ),
    .F4(\net_Lut-U117_0_S0_F_B4_to_F49_6_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S0_G_B1_to_G19_6_0 ),
    .G2(\net_cnt_lcd_reg[0]_S0_G_B2_to_G29_6_0 ),
    .G3(\net_cnt_lcd_reg[2]_S0_G_B3_to_G39_6_0 ),
    .G4(\net_cnt_lcd_reg[3]_S0_G_B4_to_G49_6_0 ),
    .XQ(),
    .X(\net_Lut-U115_1_X_to_S0_X9_6_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U144_0_0_Y_to_S0_Y9_6_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__10___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*~A2)*A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)";
  defparam iSlice__10___inst.fxmux.CONF = "F";
  defparam iSlice__10___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*~A1)";
  defparam iSlice__10___inst.gymux.CONF = "G";
  defparam iSlice__10___inst.xused.CONF = "0";
  defparam iSlice__10___inst.yused.CONF = "0";
  defparam iSlice__10___inst.f.INIT = 16'hae0c;
  defparam iSlice__10___inst.g.INIT = 16'hd000;
  SLICE iSlice__10___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U225_0_S1_F_B1_to_F19_7_0 ),
    .F2(\net_Lut-U205_0_0_S1_F_B2_to_F29_7_0 ),
    .F3(\net_Lut-U166_0_S1_F_B3_to_F39_7_0 ),
    .F4(\net_Lut-U219_0_1_S1_F_B4_to_F49_7_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[5]_S1_G_B1_to_G19_7_0 ),
    .G2(\net_cnt_lcd_reg[1]_S1_G_B2_to_G29_7_0 ),
    .G3(\net_cnt_lcd_reg[4]_S1_G_B3_to_G39_7_0 ),
    .G4(\net_Lut-U201_0_0_S1_G_B4_to_G49_7_0 ),
    .XQ(),
    .X(\net_Lut-U165_2_X_to_S1_X9_7_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U115_0_0_Y_to_S1_Y9_7_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__11___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)";
  defparam iSlice__11___inst.fxmux.CONF = "F";
  defparam iSlice__11___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*~A1)";
  defparam iSlice__11___inst.gymux.CONF = "G";
  defparam iSlice__11___inst.xused.CONF = "0";
  defparam iSlice__11___inst.yused.CONF = "0";
  defparam iSlice__11___inst.f.INIT = 16'hfefc;
  defparam iSlice__11___inst.g.INIT = 16'h4000;
  SLICE iSlice__11___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U232_0_0_S1_F_B1_to_F17_8_0 ),
    .F2(\net_Lut-U176_0_1_S1_F_B2_to_F27_8_0 ),
    .F3(\net_Lut-U175_0_0_S1_F_B3_to_F37_8_0 ),
    .F4(\net_Lut-U204_0_1_S1_F_B4_to_F47_8_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[5]_S1_G_B1_to_G17_8_0 ),
    .G2(\net_cnt_lcd_reg[3]_S1_G_B2_to_G27_8_0 ),
    .G3(\net_cnt_lcd_reg[4]_S1_G_B3_to_G37_8_0 ),
    .G4(\net_Lut-U201_0_0_S1_G_B4_to_G47_8_0 ),
    .XQ(),
    .X(\net_Lut-U174_0_X_to_S1_X7_8_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U126_0_0_Y_to_S1_Y7_8_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__12___inst.f.CONF = "#LUT:D=(((A4*~A3)*~A2)*A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__12___inst.fxmux.CONF = "F";
  defparam iSlice__12___inst.g.CONF = "#LUT:D=(((A4*~A3)*A2)*~A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__12___inst.gymux.CONF = "G";
  defparam iSlice__12___inst.xused.CONF = "0";
  defparam iSlice__12___inst.yused.CONF = "0";
  defparam iSlice__12___inst.f.INIT = 16'h307;
  defparam iSlice__12___inst.g.INIT = 16'h415;
  SLICE iSlice__12___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[7]_S0_F_B1_to_F111_9_0 ),
    .F2(\net_Lut-U232_0_0_S0_F_B2_to_F211_9_0 ),
    .F3(\net_Lut-U202_0_0_S0_F_B3_to_F311_9_0 ),
    .F4(\net_cnt_lcd_reg[2]_S0_F_B4_to_F411_9_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U230_0_0_S0_G_B1_to_G111_9_0 ),
    .G2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G211_9_0 ),
    .G3(\net_cnt_lcd_reg[5]_S0_G_B3_to_G311_9_0 ),
    .G4(\net_Lut-U198_0_0_S0_G_B4_to_G411_9_0 ),
    .XQ(),
    .X(\net_Lut-U196_4_1_X_to_S0_X11_9_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U196_5_1_Y_to_S0_Y11_9_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__13___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)";
  defparam iSlice__13___inst.fxmux.CONF = "F";
  defparam iSlice__13___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__13___inst.gymux.CONF = "G";
  defparam iSlice__13___inst.xused.CONF = "0";
  defparam iSlice__13___inst.yused.CONF = "0";
  defparam iSlice__13___inst.f.INIT = 16'h8000;
  defparam iSlice__13___inst.g.INIT = 16'h8901;
  SLICE iSlice__13___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U144_0_0_S0_F_B1_to_F18_7_0 ),
    .F2(\net_cnt_lcd_reg[4]_S0_F_B2_to_F28_7_0 ),
    .F3(\net_cnt_lcd_reg[5]_S0_F_B3_to_F38_7_0 ),
    .F4(\net_cnt_lcd_reg[6]_S0_F_B4_to_F48_7_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[3]_S0_G_B1_to_G18_7_0 ),
    .G2(\net_cnt_lcd_reg[2]_S0_G_B2_to_G28_7_0 ),
    .G3(\net_Lut-U193_0_0_S0_G_B3_to_G38_7_0 ),
    .G4(\net_Lut-U213_0_0_S0_G_B4_to_G48_7_0 ),
    .XQ(),
    .X(\net_Lut-U137_0_0_X_to_S0_X8_7_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U191_1_Y_to_S0_Y8_7_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__14___inst.f.CONF = "#LUT:D=(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__14___inst.fxmux.CONF = "F";
  defparam iSlice__14___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*A1)";
  defparam iSlice__14___inst.gymux.CONF = "G";
  defparam iSlice__14___inst.xused.CONF = "0";
  defparam iSlice__14___inst.yused.CONF = "0";
  defparam iSlice__14___inst.f.INIT = 16'h51;
  defparam iSlice__14___inst.g.INIT = 16'hddd6;
  SLICE iSlice__14___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U123_0_0_S1_F_B1_to_F110_6_0 ),
    .F2(\net_cnt_lcd_reg[5]_S1_F_B2_to_F210_6_0 ),
    .F3(\net_Lut-U124_0_0_S1_F_B3_to_F310_6_0 ),
    .F4(\net_Lut-U123_2_0_S1_F_B4_to_F410_6_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G110_6_0 ),
    .G2(\net_cnt_lcd_reg[3]_S1_G_B2_to_G210_6_0 ),
    .G3(\net_cnt_lcd_reg[2]_S1_G_B3_to_G310_6_0 ),
    .G4(\net_cnt_lcd_reg[4]_S1_G_B4_to_G410_6_0 ),
    .XQ(),
    .X(\net_Lut-U123_1_X_to_S1_X10_6_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U118_0_0_Y_to_S1_Y10_6_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__15___inst.f.CONF = "#LUT:D=(((A4*~A3)*A2)*A1)";
  defparam iSlice__15___inst.fxmux.CONF = "F";
  defparam iSlice__15___inst.g.CONF = "#LUT:D=(((A4*~A3)*~A2)*A1)";
  defparam iSlice__15___inst.gymux.CONF = "G";
  defparam iSlice__15___inst.xused.CONF = "0";
  defparam iSlice__15___inst.yused.CONF = "0";
  defparam iSlice__15___inst.f.INIT = 16'h800;
  defparam iSlice__15___inst.g.INIT = 16'h200;
  SLICE iSlice__15___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U176_0_0_S0_F_B1_to_F18_9_0 ),
    .F2(\net_cnt_lcd_reg[7]_S0_F_B2_to_F28_9_0 ),
    .F3(\net_cnt_lcd_reg[6]_S0_F_B3_to_F38_9_0 ),
    .F4(\net_cnt_lcd_reg[0]_S0_F_B4_to_F48_9_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S0_G_B1_to_G18_9_0 ),
    .G2(\net_cnt_lcd_reg[4]_S0_G_B2_to_G28_9_0 ),
    .G3(\net_cnt_lcd_reg[5]_S0_G_B3_to_G38_9_0 ),
    .G4(\net_cnt_lcd_reg[3]_S0_G_B4_to_G48_9_0 ),
    .XQ(),
    .X(\net_Lut-U176_0_1_X_to_S0_X8_9_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U204_0_1_Y_to_S0_Y8_9_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__16___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*~A2)*A1)";
  defparam iSlice__16___inst.fxmux.CONF = "F";
  defparam iSlice__16___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)";
  defparam iSlice__16___inst.gymux.CONF = "G";
  defparam iSlice__16___inst.xused.CONF = "0";
  defparam iSlice__16___inst.yused.CONF = "0";
  defparam iSlice__16___inst.f.INIT = 16'hca00;
  defparam iSlice__16___inst.g.INIT = 16'hfefc;
  SLICE iSlice__16___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U161_0_0_S0_F_B1_to_F110_8_0 ),
    .F2(\net_Lut-U215_0_0_S0_F_B2_to_F210_8_0 ),
    .F3(\net_cnt_lcd_reg[4]_S0_F_B3_to_F310_8_0 ),
    .F4(\net_Lut-U230_0_0_S0_F_B4_to_F410_8_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U205_0_0_S0_G_B1_to_G110_8_0 ),
    .G2(\net_Lut-U164_0_0_S0_G_B2_to_G210_8_0 ),
    .G3(\net_Lut-U159_0_0_S0_G_B3_to_G310_8_0 ),
    .G4(\net_Lut-U230_0_0_S0_G_B4_to_G410_8_0 ),
    .XQ(),
    .X(\net_Lut-U160_0_X_to_S0_X10_8_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U158_0_Y_to_S0_Y10_8_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__17___inst.f.CONF = "#LUT:D=(((A4*~A3)*A2)*~A1)";
  defparam iSlice__17___inst.fxmux.CONF = "F";
  defparam iSlice__17___inst.g.CONF = "#LUT:D=(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*~A1)";
  defparam iSlice__17___inst.gymux.CONF = "G";
  defparam iSlice__17___inst.xused.CONF = "0";
  defparam iSlice__17___inst.yused.CONF = "0";
  defparam iSlice__17___inst.f.INIT = 16'h400;
  defparam iSlice__17___inst.g.INIT = 16'h3074;
  SLICE iSlice__17___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[4]_S1_F_B1_to_F17_10_0 ),
    .F2(\net_cnt_lcd_reg[7]_S1_F_B2_to_F27_10_0 ),
    .F3(\net_cnt_lcd_reg[6]_S1_F_B3_to_F37_10_0 ),
    .F4(\net_cnt_lcd_reg[0]_S1_F_B4_to_F47_10_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U177_0_0_S1_G_B1_to_G17_10_0 ),
    .G2(\net_cnt_lcd_reg[4]_S1_G_B2_to_G27_10_0 ),
    .G3(\net_Lut-U129_0_S1_G_B3_to_G37_10_0 ),
    .G4(\net_Lut-U183_0_0_S1_G_B4_to_G47_10_0 ),
    .XQ(),
    .X(\net_Lut-U229_0_X_to_S1_X7_10_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U127_0_0_Y_to_S1_Y7_10_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__18___inst.f.CONF = "#LUT:D=(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__18___inst.fxmux.CONF = "F";
  defparam iSlice__18___inst.g.CONF = "#LUT:D=(((~A4*A3)*A2)*~A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__18___inst.gymux.CONF = "G";
  defparam iSlice__18___inst.xused.CONF = "0";
  defparam iSlice__18___inst.yused.CONF = "0";
  defparam iSlice__18___inst.f.INIT = 16'h3377;
  defparam iSlice__18___inst.g.INIT = 16'h45;
  SLICE iSlice__18___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[7]_S0_F_B1_to_F110_7_0 ),
    .F2(\net_Lut-U232_0_0_S0_F_B2_to_F210_7_0 ),
    .F3(\net_cnt_lcd_reg[4]_S0_F_B3_to_F310_7_0 ),
    .F4(\net_cnt_lcd_reg[2]_S0_F_B4_to_F410_7_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U230_0_0_S0_G_B1_to_G110_7_0 ),
    .G2(\net_cnt_lcd_reg[4]_S0_G_B2_to_G210_7_0 ),
    .G3(\net_Lut-U201_0_0_S0_G_B3_to_G310_7_0 ),
    .G4(\net_Lut-U197_0_0_S0_G_B4_to_G410_7_0 ),
    .XQ(),
    .X(\net_Lut-U196_6_1_X_to_S0_X10_7_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U196_7_1_Y_to_S0_Y10_7_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__19___inst.f.CONF = "#LUT:D=(((~A4*~A3)*A2)*~A1)";
  defparam iSlice__19___inst.fxmux.CONF = "F";
  defparam iSlice__19___inst.g.CONF = "#LUT:D=(((A4*~A3)*~A2)*~A1)";
  defparam iSlice__19___inst.gymux.CONF = "G";
  defparam iSlice__19___inst.xused.CONF = "0";
  defparam iSlice__19___inst.yused.CONF = "0";
  defparam iSlice__19___inst.f.INIT = 16'h4;
  defparam iSlice__19___inst.g.INIT = 16'h100;
  SLICE iSlice__19___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[5]_S0_F_B1_to_F110_10_0 ),
    .F2(\net_cnt_lcd_reg[4]_S0_F_B2_to_F210_10_0 ),
    .F3(\net_cnt_lcd_reg[2]_S0_F_B3_to_F310_10_0 ),
    .F4(\net_cnt_lcd_reg[3]_S0_F_B4_to_F410_10_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[4]_S0_G_B1_to_G110_10_0 ),
    .G2(\net_cnt_lcd_reg[7]_S0_G_B2_to_G210_10_0 ),
    .G3(\net_cnt_lcd_reg[6]_S0_G_B3_to_G310_10_0 ),
    .G4(\net_cnt_lcd_reg[0]_S0_G_B4_to_G410_10_0 ),
    .XQ(),
    .X(\net_Lut-U217_1_X_to_S0_X10_10_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U224_0_0_Y_to_S0_Y10_10_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__20___inst.f.CONF = "#LUT:D=(((A4*~A3)*~A2)*A1)";
  defparam iSlice__20___inst.fxmux.CONF = "F";
  defparam iSlice__20___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*~A2)*A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*~A3)*A2)*A1)";
  defparam iSlice__20___inst.gymux.CONF = "G";
  defparam iSlice__20___inst.xused.CONF = "0";
  defparam iSlice__20___inst.yused.CONF = "0";
  defparam iSlice__20___inst.f.INIT = 16'h200;
  defparam iSlice__20___inst.g.INIT = 16'h6b08;
  SLICE iSlice__20___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[2]_S0_F_B1_to_F17_9_0 ),
    .F2(\net_cnt_lcd_reg[7]_S0_F_B2_to_F27_9_0 ),
    .F3(\net_cnt_lcd_reg[6]_S0_F_B3_to_F37_9_0 ),
    .F4(\net_cnt_lcd_reg[0]_S0_F_B4_to_F47_9_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[2]_S0_G_B1_to_G17_9_0 ),
    .G2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G27_9_0 ),
    .G3(\net_cnt_lcd_reg[5]_S0_G_B3_to_G37_9_0 ),
    .G4(\net_cnt_lcd_reg[3]_S0_G_B4_to_G47_9_0 ),
    .XQ(),
    .X(\net_Lut-U201_0_0_X_to_S0_X7_9_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U132_0_Y_to_S0_Y7_9_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__21___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*~A2)*A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__21___inst.fxmux.CONF = "F";
  defparam iSlice__21___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__21___inst.gymux.CONF = "G";
  defparam iSlice__21___inst.xused.CONF = "0";
  defparam iSlice__21___inst.yused.CONF = "0";
  defparam iSlice__21___inst.f.INIT = 16'hf73b;
  defparam iSlice__21___inst.g.INIT = 16'hf755;
  SLICE iSlice__21___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[4]_S1_F_B1_to_F19_6_0 ),
    .F2(\net_Lut-U232_0_0_S1_F_B2_to_F29_6_0 ),
    .F3(\net_cnt_lcd_reg[7]_S1_F_B3_to_F39_6_0 ),
    .F4(\net_cnt_lcd_reg[5]_S1_F_B4_to_F49_6_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G19_6_0 ),
    .G2(\net_cnt_lcd_reg[5]_S1_G_B2_to_G29_6_0 ),
    .G3(\net_cnt_lcd_reg[2]_S1_G_B3_to_G39_6_0 ),
    .G4(\net_cnt_lcd_reg[3]_S1_G_B4_to_G49_6_0 ),
    .XQ(),
    .X(\net_Lut-U166_0_X_to_S1_X9_6_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U122_0_0_Y_to_S1_Y9_6_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__22___inst.f.CONF = "#LUT:D=((~A3*A2)*~A1)+((~A3*~A2)*A1)+((~A3*~A2)*~A1)";
  defparam iSlice__22___inst.fxmux.CONF = "F";
  defparam iSlice__22___inst.g.CONF = "#LUT:D=((~A3*~A2)*~A1)";
  defparam iSlice__22___inst.gymux.CONF = "G";
  defparam iSlice__22___inst.xused.CONF = "0";
  defparam iSlice__22___inst.yused.CONF = "0";
  defparam iSlice__22___inst.f.INIT = 16'h7;
  defparam iSlice__22___inst.g.INIT = 16'h1;
  SLICE iSlice__22___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U153_0_S1_F_B1_to_F19_8_0 ),
    .F2(\net_Lut-U225_0_S1_F_B2_to_F29_8_0 ),
    .F3(\net_Lut-U151_0_S1_F_B3_to_F39_8_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U162_0_0_S1_G_B1_to_G19_8_0 ),
    .G2(\net_Lut-U165_2_S1_G_B2_to_G29_8_0 ),
    .G3(\net_Lut-U164_0_0_S1_G_B3_to_G39_8_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U150_0_X_to_S1_X9_8_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U162_1_Y_to_S1_Y9_8_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__23___inst.f.CONF = "#LUT:D=((A3*A2)*A1)+((A3*~A2)*~A1)+((~A3*A2)*~A1)+((~A3*~A2)*~A1)";
  defparam iSlice__23___inst.fxmux.CONF = "F";
  defparam iSlice__23___inst.g.CONF = "#LUT:D=((~A3*~A2)*~A1)";
  defparam iSlice__23___inst.gymux.CONF = "G";
  defparam iSlice__23___inst.xused.CONF = "0";
  defparam iSlice__23___inst.yused.CONF = "0";
  defparam iSlice__23___inst.f.INIT = 16'h95;
  defparam iSlice__23___inst.g.INIT = 16'h1;
  SLICE iSlice__23___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[5]_S1_F_B1_to_F17_7_0 ),
    .F2(\net_Lut-U144_0_0_S1_F_B2_to_F27_7_0 ),
    .F3(\net_cnt_lcd_reg[4]_S1_F_B3_to_F37_7_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U191_1_S1_G_B1_to_G17_7_0 ),
    .G2(\net_Lut-U178_0_S1_G_B2_to_G27_7_0 ),
    .G3(\net_Lut-U174_0_S1_G_B3_to_G37_7_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U141_0_X_to_S1_X7_7_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U173_1_Y_to_S1_Y7_7_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__24___inst.f.CONF = "#LUT:D=((A3*~A2)*~A1)";
  defparam iSlice__24___inst.fxmux.CONF = "F";
  defparam iSlice__24___inst.g.CONF = "#LUT:D=((~A3*A2)*A1)+((~A3*~A2)*A1)+((~A3*~A2)*~A1)";
  defparam iSlice__24___inst.gymux.CONF = "G";
  defparam iSlice__24___inst.xused.CONF = "0";
  defparam iSlice__24___inst.yused.CONF = "0";
  defparam iSlice__24___inst.f.INIT = 16'h10;
  defparam iSlice__24___inst.g.INIT = 16'hb;
  SLICE iSlice__24___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[7]_S1_F_B1_to_F110_10_0 ),
    .F2(\net_cnt_lcd_reg[6]_S1_F_B2_to_F210_10_0 ),
    .F3(\net_cnt_lcd_reg[0]_S1_F_B3_to_F310_10_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[2]_S1_G_B1_to_G110_10_0 ),
    .G2(\net_Lut-U223_0_S1_G_B2_to_G210_10_0 ),
    .G3(\net_Lut-U208_0_S1_G_B3_to_G310_10_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U225_0_X_to_S1_X10_10_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U195_0_Y_to_S1_Y10_10_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__25___inst.f.CONF = "#LUT:D=((A3*A2)*~A1)+((A3*~A2)*~A1)+((~A3*A2)*~A1)";
  defparam iSlice__25___inst.fxmux.CONF = "F";
  defparam iSlice__25___inst.g.CONF = "#LUT:D=((A3*~A2)*A1)";
  defparam iSlice__25___inst.gymux.CONF = "G";
  defparam iSlice__25___inst.xused.CONF = "0";
  defparam iSlice__25___inst.yused.CONF = "0";
  defparam iSlice__25___inst.f.INIT = 16'h54;
  defparam iSlice__25___inst.g.INIT = 16'h20;
  SLICE iSlice__25___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[1]_S0_F_B1_to_F19_8_0 ),
    .F2(\net_Lut-U170_1_S0_F_B2_to_F29_8_0 ),
    .F3(\net_Lut-U224_0_1_S0_F_B3_to_F39_8_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U190_0_1_S0_G_B1_to_G19_8_0 ),
    .G2(\net_cnt_lcd_reg[4]_S0_G_B2_to_G29_8_0 ),
    .G3(\net_Lut-U201_0_0_S0_G_B3_to_G39_8_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U162_0_0_X_to_S0_X9_8_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U164_0_0_Y_to_S0_Y9_8_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__26___inst.f.CONF = "#LUT:D=(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__26___inst.fxmux.CONF = "F";
  defparam iSlice__26___inst.g.CONF = "#LUT:D=(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__26___inst.gymux.CONF = "G";
  defparam iSlice__26___inst.xused.CONF = "0";
  defparam iSlice__26___inst.yused.CONF = "0";
  defparam iSlice__26___inst.f.INIT = 16'h1;
  defparam iSlice__26___inst.g.INIT = 16'h111;
  SLICE iSlice__26___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U205_0_0_S0_F_B1_to_F111_8_0 ),
    .F2(\net_Lut-U204_0_1_S0_F_B2_to_F211_8_0 ),
    .F3(\net_Lut-U202_0_0_S0_F_B3_to_F311_8_0 ),
    .F4(\net_Lut-U201_0_0_S0_F_B4_to_F411_8_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U205_0_0_S0_G_B1_to_G111_8_0 ),
    .G2(\net_Lut-U204_0_1_S0_G_B2_to_G211_8_0 ),
    .G3(\net_cnt_lcd_reg[1]_S0_G_B3_to_G311_8_0 ),
    .G4(\net_cnt_lcd_reg[5]_S0_G_B4_to_G411_8_0 ),
    .XQ(),
    .X(\net_Lut-U196_0_1_X_to_S0_X11_8_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U196_1_0_Y_to_S0_Y11_8_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__27___inst.f.CONF = "#LUT:D=((A3*A2)*A1)+((A3*A2)*~A1)+((A3*~A2)*A1)+((~A3*~A2)*A1)";
  defparam iSlice__27___inst.fxmux.CONF = "F";
  defparam iSlice__27___inst.g.CONF = "#LUT:D=((~A3*~A2)*A1)";
  defparam iSlice__27___inst.gymux.CONF = "G";
  defparam iSlice__27___inst.xused.CONF = "0";
  defparam iSlice__27___inst.yused.CONF = "0";
  defparam iSlice__27___inst.f.INIT = 16'he2;
  defparam iSlice__27___inst.g.INIT = 16'h2;
  SLICE iSlice__27___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U189_2_S0_F_B1_to_F18_8_0 ),
    .F2(\net_cnt_lcd_reg[4]_S0_F_B2_to_F28_8_0 ),
    .F3(\net_Lut-U179_2_S0_F_B3_to_F38_8_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U213_0_0_S0_G_B1_to_G18_8_0 ),
    .G2(\net_cnt_lcd_reg[2]_S0_G_B2_to_G28_8_0 ),
    .G3(\net_cnt_lcd_reg[3]_S0_G_B3_to_G38_8_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U178_0_X_to_S0_X8_8_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U209_0_0_Y_to_S0_Y8_8_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__28___inst.f.CONF = "#LUT:D=((A3*A2)*A1)+((A3*~A2)*A1)+((~A3*~A2)*A1)";
  defparam iSlice__28___inst.fxmux.CONF = "F";
  defparam iSlice__28___inst.g.CONF = "#LUT:D=((A3*~A2)*A1)";
  defparam iSlice__28___inst.gymux.CONF = "G";
  defparam iSlice__28___inst.xused.CONF = "0";
  defparam iSlice__28___inst.yused.CONF = "0";
  defparam iSlice__28___inst.f.INIT = 16'ha2;
  defparam iSlice__28___inst.g.INIT = 16'h20;
  SLICE iSlice__28___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U154_0_S0_F_B1_to_F19_9_0 ),
    .F2(\net_cnt_lcd_reg[4]_S0_F_B2_to_F29_9_0 ),
    .F3(\net_cnt_lcd_reg[3]_S0_F_B3_to_F39_9_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[7]_S0_G_B1_to_G19_9_0 ),
    .G2(\net_cnt_lcd_reg[6]_S0_G_B2_to_G29_9_0 ),
    .G3(\net_cnt_lcd_reg[0]_S0_G_B3_to_G39_9_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U154_1_X_to_S0_X9_9_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U230_0_0_Y_to_S0_Y9_9_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__29___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*A2)*A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__29___inst.fxmux.CONF = "F";
  defparam iSlice__29___inst.g.CONF = "#LUT:D=(((A4*~A3)*A2)*A1)";
  defparam iSlice__29___inst.gymux.CONF = "G";
  defparam iSlice__29___inst.xused.CONF = "0";
  defparam iSlice__29___inst.yused.CONF = "0";
  defparam iSlice__29___inst.f.INIT = 16'hbf8f;
  defparam iSlice__29___inst.g.INIT = 16'h800;
  SLICE iSlice__29___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[4]_S1_F_B1_to_F18_7_0 ),
    .F2(\net_cnt_lcd_reg[7]_S1_F_B2_to_F28_7_0 ),
    .F3(\net_Lut-U232_0_0_S1_F_B3_to_F38_7_0 ),
    .F4(\net_cnt_lcd_reg[5]_S1_F_B4_to_F48_7_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[4]_S1_G_B1_to_G18_7_0 ),
    .G2(\net_cnt_lcd_reg[7]_S1_G_B2_to_G28_7_0 ),
    .G3(\net_cnt_lcd_reg[6]_S1_G_B3_to_G38_7_0 ),
    .G4(\net_cnt_lcd_reg[0]_S1_G_B4_to_G48_7_0 ),
    .XQ(),
    .X(\net_Lut-U193_0_0_X_to_S1_X8_7_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U213_0_0_Y_to_S1_Y8_7_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__30___inst.ckinv.CONF = "1";
  defparam iSlice__30___inst.dxmux.CONF = "1";
  defparam iSlice__30___inst.dymux.CONF = "1";
  defparam iSlice__30___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__30___inst.ffx.TYPE = "#FF";
  defparam iSlice__30___inst.ffy.TYPE = "#FF";
  defparam iSlice__30___inst.fxmux.CONF = "F";
  defparam iSlice__30___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__30___inst.gymux.CONF = "G";
  defparam iSlice__30___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__30___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__30___inst.srffmux.CONF = "0";
  defparam iSlice__30___inst.srmux.CONF = "SR_B";
  defparam iSlice__30___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__30___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__30___inst.f.INIT = 16'h5;
  defparam iSlice__30___inst.g.INIT = 16'h5;
  SLICE iSlice__30___inst (
    .CIN(),
    .SR(net_rst_nInvLut_S0_SR_B_to_SR7_3_0),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK7_3_0 ),
    .CE(),
    .BX(),
    .F1(\net_Lut-U173_1_S0_F_B1_to_F17_3_0 ),
    .F2(net_U113_S0_F_B2_to_F27_3_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U126_1_S0_G_B1_to_G17_3_0 ),
    .G2(net_U113_S0_G_B2_to_G27_3_0),
    .G3(),
    .G4(),
    .XQ(\net_lcd_db_reg[3]_XQ_to_S0_XQ7_3_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_lcd_db_reg[0]_YQ_to_S0_YQ7_3_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__31___inst.ckinv.CONF = "1";
  defparam iSlice__31___inst.dxmux.CONF = "1";
  defparam iSlice__31___inst.dymux.CONF = "1";
  defparam iSlice__31___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__31___inst.ffx.TYPE = "#FF";
  defparam iSlice__31___inst.ffy.TYPE = "#FF";
  defparam iSlice__31___inst.fxmux.CONF = "F";
  defparam iSlice__31___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__31___inst.gymux.CONF = "G";
  defparam iSlice__31___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__31___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__31___inst.srffmux.CONF = "0";
  defparam iSlice__31___inst.srmux.CONF = "SR_B";
  defparam iSlice__31___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__31___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__31___inst.f.INIT = 16'h5;
  defparam iSlice__31___inst.g.INIT = 16'h5;
  SLICE iSlice__31___inst (
    .CIN(),
    .SR(net_rst_nInvLut_S0_SR_B_to_SR9_3_0),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK9_3_0 ),
    .CE(),
    .BX(),
    .F1(\net_Lut-U150_0_S0_F_B1_to_F19_3_0 ),
    .F2(net_U113_S0_F_B2_to_F29_3_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U157_1_S0_G_B1_to_G19_3_0 ),
    .G2(net_U113_S0_G_B2_to_G29_3_0),
    .G3(),
    .G4(),
    .XQ(\net_lcd_db_reg[6]_XQ_to_S0_XQ9_3_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_lcd_db_reg[5]_YQ_to_S0_YQ9_3_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__32___inst.ckinv.CONF = "1";
  defparam iSlice__32___inst.dxmux.CONF = "1";
  defparam iSlice__32___inst.dymux.CONF = "1";
  defparam iSlice__32___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__32___inst.ffx.TYPE = "#FF";
  defparam iSlice__32___inst.ffy.TYPE = "#FF";
  defparam iSlice__32___inst.fxmux.CONF = "F";
  defparam iSlice__32___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__32___inst.gymux.CONF = "G";
  defparam iSlice__32___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__32___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__32___inst.srffmux.CONF = "0";
  defparam iSlice__32___inst.srmux.CONF = "SR_B";
  defparam iSlice__32___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__32___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__32___inst.f.INIT = 16'h5;
  defparam iSlice__32___inst.g.INIT = 16'h5;
  SLICE iSlice__32___inst (
    .CIN(),
    .SR(net_rst_nInvLut_S0_SR_B_to_SR9_4_0),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK9_4_0 ),
    .CE(),
    .BX(),
    .F1(\net_Lut-U195_1_S0_F_B1_to_F19_4_0 ),
    .F2(net_U113_S0_F_B2_to_F29_4_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U162_1_S0_G_B1_to_G19_4_0 ),
    .G2(net_U113_S0_G_B2_to_G29_4_0),
    .G3(),
    .G4(),
    .XQ(\net_lcd_db_reg[2]_XQ_to_S0_XQ9_4_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_lcd_db_reg[4]_YQ_to_S0_YQ9_4_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__33___inst.ckinv.CONF = "1";
  defparam iSlice__33___inst.dxmux.CONF = "1";
  defparam iSlice__33___inst.dymux.CONF = "1";
  defparam iSlice__33___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__33___inst.ffx.TYPE = "#FF";
  defparam iSlice__33___inst.ffy.TYPE = "#FF";
  defparam iSlice__33___inst.fxmux.CONF = "F";
  defparam iSlice__33___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__33___inst.gymux.CONF = "G";
  defparam iSlice__33___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__33___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__33___inst.srffmux.CONF = "0";
  defparam iSlice__33___inst.srmux.CONF = "SR_B";
  defparam iSlice__33___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__33___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__33___inst.f.INIT = 16'h5;
  defparam iSlice__33___inst.g.INIT = 16'h5;
  SLICE iSlice__33___inst (
    .CIN(),
    .SR(net_rst_nInvLut_S1_SR_B_to_SR7_6_0),
    .CLK(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK7_6_0 ),
    .CE(),
    .BX(),
    .F1(\net_Lut-U138_0_S1_F_B1_to_F17_6_0 ),
    .F2(net_U113_S1_F_B2_to_F27_6_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U136_0_S1_G_B1_to_G17_6_0 ),
    .G2(net_U113_S1_G_B2_to_G27_6_0),
    .G3(),
    .G4(),
    .XQ(\net_cnt_lcd_reg[6]_XQ_to_S1_XQ7_6_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_cnt_lcd_reg[7]_YQ_to_S1_YQ7_6_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__34___inst.f.CONF = "#LUT:D=(((A4*A3)*~A2)*A1)";
  defparam iSlice__34___inst.fxmux.CONF = "F";
  defparam iSlice__34___inst.g.CONF = "#LUT:D=(((A4*A3)*~A2)*A1)";
  defparam iSlice__34___inst.gymux.CONF = "G";
  defparam iSlice__34___inst.xused.CONF = "0";
  defparam iSlice__34___inst.yused.CONF = "0";
  defparam iSlice__34___inst.f.INIT = 16'h2000;
  defparam iSlice__34___inst.g.INIT = 16'h2000;
  SLICE iSlice__34___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[7]_S0_F_B1_to_F110_9_0 ),
    .F2(\net_cnt_lcd_reg[6]_S0_F_B2_to_F210_9_0 ),
    .F3(\net_cnt_lcd_reg[0]_S0_F_B3_to_F310_9_0 ),
    .F4(\net_Lut-U217_1_S0_F_B4_to_F410_9_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[7]_S0_G_B1_to_G110_9_0 ),
    .G2(\net_cnt_lcd_reg[6]_S0_G_B2_to_G210_9_0 ),
    .G3(\net_cnt_lcd_reg[0]_S0_G_B3_to_G310_9_0 ),
    .G4(\net_cnt_lcd_reg[5]_S0_G_B4_to_G410_9_0 ),
    .XQ(),
    .X(\net_Lut-U152_0_0_X_to_S0_X10_9_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U170_0_Y_to_S0_Y10_9_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__35___inst.ckinv.CONF = "1";
  defparam iSlice__35___inst.dxmux.CONF = "1";
  defparam iSlice__35___inst.dymux.CONF = "1";
  defparam iSlice__35___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__35___inst.ffx.TYPE = "#FF";
  defparam iSlice__35___inst.ffy.TYPE = "#FF";
  defparam iSlice__35___inst.fxmux.CONF = "F";
  defparam iSlice__35___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__35___inst.gymux.CONF = "G";
  defparam iSlice__35___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__35___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__35___inst.srffmux.CONF = "0";
  defparam iSlice__35___inst.srmux.CONF = "SR_B";
  defparam iSlice__35___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__35___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__35___inst.f.INIT = 16'h5;
  defparam iSlice__35___inst.g.INIT = 16'h5;
  SLICE iSlice__35___inst (
    .CIN(),
    .SR(net_rst_nInvLut_S0_SR_B_to_SR9_5_0),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK9_5_0 ),
    .CE(),
    .BX(),
    .F1(\net_Lut-U147_0_S0_F_B1_to_F19_5_0 ),
    .F2(net_U113_S0_F_B2_to_F29_5_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U145_0_S0_G_B1_to_G19_5_0 ),
    .G2(net_U113_S0_G_B2_to_G29_5_0),
    .G3(),
    .G4(),
    .XQ(\net_cnt_lcd_reg[2]_XQ_to_S0_XQ9_5_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_cnt_lcd_reg[3]_YQ_to_S0_YQ9_5_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__36___inst.ckinv.CONF = "1";
  defparam iSlice__36___inst.dxmux.CONF = "1";
  defparam iSlice__36___inst.dymux.CONF = "1";
  defparam iSlice__36___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__36___inst.ffx.TYPE = "#FF";
  defparam iSlice__36___inst.ffy.TYPE = "#FF";
  defparam iSlice__36___inst.fxmux.CONF = "F";
  defparam iSlice__36___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__36___inst.gymux.CONF = "G";
  defparam iSlice__36___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__36___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__36___inst.srffmux.CONF = "0";
  defparam iSlice__36___inst.srmux.CONF = "SR_B";
  defparam iSlice__36___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__36___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__36___inst.f.INIT = 16'h5;
  defparam iSlice__36___inst.g.INIT = 16'h5;
  SLICE iSlice__36___inst (
    .CIN(),
    .SR(net_rst_nInvLut_S0_SR_B_to_SR7_6_0),
    .CLK(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK7_6_0 ),
    .CE(),
    .BX(),
    .F1(\net_Lut-U143_0_S0_F_B1_to_F17_6_0 ),
    .F2(net_U113_S0_F_B2_to_F27_6_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U141_0_S0_G_B1_to_G17_6_0 ),
    .G2(net_U113_S0_G_B2_to_G27_6_0),
    .G3(),
    .G4(),
    .XQ(\net_cnt_lcd_reg[4]_XQ_to_S0_XQ7_6_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_cnt_lcd_reg[5]_YQ_to_S0_YQ7_6_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__37___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__37___inst.fxmux.CONF = "F";
  defparam iSlice__37___inst.g.CONF = "#LUT:D=((A3*A2)*A1)+((A3*~A2)*~A1)+((~A3*A2)*~A1)+((~A3*~A2)*~A1)";
  defparam iSlice__37___inst.gymux.CONF = "G";
  defparam iSlice__37___inst.xused.CONF = "0";
  defparam iSlice__37___inst.yused.CONF = "0";
  defparam iSlice__37___inst.f.INIT = 16'h5;
  defparam iSlice__37___inst.g.INIT = 16'h95;
  SLICE iSlice__37___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Buf-pad-rst_n_S1_F_B1_to_F19_5_0 ),
    .F2(net_U113_S1_F_B2_to_F29_5_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[2]_S1_G_B1_to_G19_5_0 ),
    .G2(\net_cnt_lcd_reg[1]_S1_G_B2_to_G29_5_0 ),
    .G3(\net_cnt_lcd_reg[0]_S1_G_B3_to_G39_5_0 ),
    .G4(),
    .XQ(),
    .X(net_rst_nInvLut_X_to_S1_X9_5_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U147_0_Y_to_S1_Y9_5_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__38___inst.f.CONF = "#LUT:D=((~A3*A2)*~A1)";
  defparam iSlice__38___inst.fxmux.CONF = "F";
  defparam iSlice__38___inst.g.CONF = "#LUT:D=((~A3*~A2)*A1)";
  defparam iSlice__38___inst.gymux.CONF = "G";
  defparam iSlice__38___inst.xused.CONF = "0";
  defparam iSlice__38___inst.yused.CONF = "0";
  defparam iSlice__38___inst.f.INIT = 16'h4;
  defparam iSlice__38___inst.g.INIT = 16'h2;
  SLICE iSlice__38___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[4]_S1_F_B1_to_F110_7_0 ),
    .F2(\net_Lut-U201_0_0_S1_F_B2_to_F210_7_0 ),
    .F3(\net_Lut-U182_0_1_S1_F_B3_to_F310_7_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[4]_S1_G_B1_to_G110_7_0 ),
    .G2(\net_cnt_lcd_reg[3]_S1_G_B2_to_G210_7_0 ),
    .G3(\net_cnt_lcd_reg[1]_S1_G_B3_to_G310_7_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U159_0_0_X_to_S1_X10_7_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U197_0_0_Y_to_S1_Y10_7_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__39___inst.f.CONF = "#LUT:D=((A3*A2)*~A1)+((A3*~A2)*A1)+((~A3*A2)*A1)+((~A3*A2)*~A1)+((~A3*~A2)*~A1)";
  defparam iSlice__39___inst.fxmux.CONF = "F";
  defparam iSlice__39___inst.g.CONF = "#LUT:D=((A3*~A2)*~A1)";
  defparam iSlice__39___inst.gymux.CONF = "G";
  defparam iSlice__39___inst.xused.CONF = "0";
  defparam iSlice__39___inst.yused.CONF = "0";
  defparam iSlice__39___inst.f.INIT = 16'h6d;
  defparam iSlice__39___inst.g.INIT = 16'h10;
  SLICE iSlice__39___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[1]_S0_F_B1_to_F19_7_0 ),
    .F2(\net_cnt_lcd_reg[5]_S0_F_B2_to_F29_7_0 ),
    .F3(\net_cnt_lcd_reg[3]_S0_F_B3_to_F39_7_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S0_G_B1_to_G19_7_0 ),
    .G2(\net_cnt_lcd_reg[2]_S0_G_B2_to_G29_7_0 ),
    .G3(\net_Lut-U213_0_0_S0_G_B3_to_G39_7_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U182_0_1_X_to_S0_X9_7_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U211_0_0_Y_to_S0_Y9_7_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__40___inst.f.CONF = "#LUT:D=((A3*~A2)*A1)";
  defparam iSlice__40___inst.fxmux.CONF = "F";
  defparam iSlice__40___inst.g.CONF = "#LUT:D=((A3*~A2)*A1)";
  defparam iSlice__40___inst.gymux.CONF = "G";
  defparam iSlice__40___inst.xused.CONF = "0";
  defparam iSlice__40___inst.yused.CONF = "0";
  defparam iSlice__40___inst.f.INIT = 16'h20;
  defparam iSlice__40___inst.g.INIT = 16'h20;
  SLICE iSlice__40___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U201_0_0_S0_F_B1_to_F17_7_0 ),
    .F2(\net_cnt_lcd_reg[5]_S0_F_B2_to_F27_7_0 ),
    .F3(\net_cnt_lcd_reg[3]_S0_F_B3_to_F37_7_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S0_G_B1_to_G17_7_0 ),
    .G2(\net_cnt_lcd_reg[3]_S0_G_B2_to_G27_7_0 ),
    .G3(\net_cnt_lcd_reg[2]_S0_G_B3_to_G37_7_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U175_0_0_X_to_S0_X7_7_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U205_0_0_Y_to_S0_Y7_7_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__41___inst.f.CONF = "#LUT:D=((A3*A2)*~A1)";
  defparam iSlice__41___inst.fxmux.CONF = "F";
  defparam iSlice__41___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__41___inst.gymux.CONF = "G";
  defparam iSlice__41___inst.xused.CONF = "0";
  defparam iSlice__41___inst.yused.CONF = "0";
  defparam iSlice__41___inst.f.INIT = 16'h40;
  defparam iSlice__41___inst.g.INIT = 16'h9555;
  SLICE iSlice__41___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[5]_S0_F_B1_to_F110_5_0 ),
    .F2(\net_cnt_lcd_reg[3]_S0_F_B2_to_F210_5_0 ),
    .F3(\net_cnt_lcd_reg[2]_S0_F_B3_to_F310_5_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[3]_S0_G_B1_to_G110_5_0 ),
    .G2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G210_5_0 ),
    .G3(\net_cnt_lcd_reg[0]_S0_G_B3_to_G310_5_0 ),
    .G4(\net_cnt_lcd_reg[2]_S0_G_B4_to_G410_5_0 ),
    .XQ(),
    .X(\net_Lut-U123_0_0_X_to_S0_X10_5_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U145_0_Y_to_S0_Y10_5_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__42___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__42___inst.fxmux.CONF = "F";
  defparam iSlice__42___inst.g.CONF = "#LUT:D=(((~A4*A3)*~A2)*~A1)";
  defparam iSlice__42___inst.gymux.CONF = "G";
  defparam iSlice__42___inst.xused.CONF = "0";
  defparam iSlice__42___inst.yused.CONF = "0";
  defparam iSlice__42___inst.f.INIT = 16'h6d65;
  defparam iSlice__42___inst.g.INIT = 16'h10;
  SLICE iSlice__42___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[1]_S1_F_B1_to_F18_9_0 ),
    .F2(\net_cnt_lcd_reg[5]_S1_F_B2_to_F28_9_0 ),
    .F3(\net_cnt_lcd_reg[3]_S1_F_B3_to_F38_9_0 ),
    .F4(\net_cnt_lcd_reg[2]_S1_F_B4_to_F48_9_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G18_9_0 ),
    .G2(\net_cnt_lcd_reg[5]_S1_G_B2_to_G28_9_0 ),
    .G3(\net_cnt_lcd_reg[4]_S1_G_B3_to_G38_9_0 ),
    .G4(\net_cnt_lcd_reg[2]_S1_G_B4_to_G48_9_0 ),
    .XQ(),
    .X(\net_Lut-U180_0_0_X_to_S1_X8_9_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U176_0_0_Y_to_S1_Y8_9_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__43___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*A2)*~A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)";
  defparam iSlice__43___inst.fxmux.CONF = "F";
  defparam iSlice__43___inst.g.CONF = "#LUT:D=(((A4*~A3)*~A2)*A1)";
  defparam iSlice__43___inst.gymux.CONF = "G";
  defparam iSlice__43___inst.xused.CONF = "0";
  defparam iSlice__43___inst.yused.CONF = "0";
  defparam iSlice__43___inst.f.INIT = 16'hfdcc;
  defparam iSlice__43___inst.g.INIT = 16'h200;
  SLICE iSlice__43___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[4]_S0_F_B1_to_F111_6_0 ),
    .F2(\net_cnt_lcd_reg[3]_S0_F_B2_to_F211_6_0 ),
    .F3(\net_cnt_lcd_reg[1]_S0_F_B3_to_F311_6_0 ),
    .F4(\net_cnt_lcd_reg[2]_S0_F_B4_to_F411_6_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[4]_S0_G_B1_to_G111_6_0 ),
    .G2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G211_6_0 ),
    .G3(\net_cnt_lcd_reg[5]_S0_G_B3_to_G311_6_0 ),
    .G4(\net_cnt_lcd_reg[3]_S0_G_B4_to_G411_6_0 ),
    .XQ(),
    .X(\net_Lut-U124_0_0_X_to_S0_X11_6_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U123_2_0_Y_to_S0_Y11_6_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__44___inst.f.CONF = "#LUT:D=(A2*A1)+(~A2*~A1)";
  defparam iSlice__44___inst.fxmux.CONF = "F";
  defparam iSlice__44___inst.g.CONF = "#LUT:D=(A2*A1)+(~A2*~A1)";
  defparam iSlice__44___inst.gymux.CONF = "G";
  defparam iSlice__44___inst.xused.CONF = "0";
  defparam iSlice__44___inst.yused.CONF = "0";
  defparam iSlice__44___inst.f.INIT = 16'h9;
  defparam iSlice__44___inst.g.INIT = 16'h9;
  SLICE iSlice__44___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[4]_S0_F_B1_to_F18_6_0 ),
    .F2(\net_Lut-U144_0_0_S0_F_B2_to_F28_6_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[7]_S0_G_B1_to_G18_6_0 ),
    .G2(\net_Lut-U137_0_0_S0_G_B2_to_G28_6_0 ),
    .G3(),
    .G4(),
    .XQ(),
    .X(\net_Lut-U143_0_X_to_S0_X8_6_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U136_0_Y_to_S0_Y8_6_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__45___inst.f.CONF = "#LUT:D=(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__45___inst.fxmux.CONF = "F";
  defparam iSlice__45___inst.g.CONF = "#LUT:D=(((A4*A3)*~A2)*~A1)+(((~A4*A3)*~A2)*~A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__45___inst.gymux.CONF = "G";
  defparam iSlice__45___inst.xused.CONF = "0";
  defparam iSlice__45___inst.yused.CONF = "0";
  defparam iSlice__45___inst.f.INIT = 16'h11;
  defparam iSlice__45___inst.g.INIT = 16'h1011;
  SLICE iSlice__45___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U205_0_0_S1_F_B1_to_F111_7_0 ),
    .F2(\net_Lut-U204_0_1_S1_F_B2_to_F211_7_0 ),
    .F3(\net_cnt_lcd_reg[4]_S1_F_B3_to_F311_7_0 ),
    .F4(\net_Lut-U201_0_0_S1_F_B4_to_F411_7_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U205_0_0_S1_G_B1_to_G111_7_0 ),
    .G2(\net_Lut-U204_0_1_S1_G_B2_to_G211_7_0 ),
    .G3(\net_cnt_lcd_reg[4]_S1_G_B3_to_G311_7_0 ),
    .G4(\net_Lut-U201_0_0_S1_G_B4_to_G411_7_0 ),
    .XQ(),
    .X(\net_Lut-U196_2_1_X_to_S1_X11_7_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U196_3_0_Y_to_S1_Y11_7_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__46___inst.f.CONF = "#LUT:D=(~A2*~A1)";
  defparam iSlice__46___inst.fxmux.CONF = "F";
  defparam iSlice__46___inst.g.CONF = "#LUT:D=(~A2*A1)";
  defparam iSlice__46___inst.gymux.CONF = "G";
  defparam iSlice__46___inst.xused.CONF = "0";
  defparam iSlice__46___inst.yused.CONF = "0";
  defparam iSlice__46___inst.f.INIT = 16'h1;
  defparam iSlice__46___inst.g.INIT = 16'h2;
  SLICE iSlice__46___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U216_0_0_S0_F_B1_to_F111_10_0 ),
    .F2(\net_Lut-U217_1_S0_F_B2_to_F211_10_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[4]_S0_G_B1_to_G111_10_0 ),
    .G2(\net_cnt_lcd_reg[3]_S0_G_B2_to_G211_10_0 ),
    .G3(),
    .G4(),
    .XQ(),
    .X(\net_Lut-U216_0_X_to_S0_X11_10_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U198_0_0_Y_to_S0_Y11_10_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__47___inst.ckinv.CONF = "1";
  defparam iSlice__47___inst.dxmux.CONF = "1";
  defparam iSlice__47___inst.dymux.CONF = "1";
  defparam iSlice__47___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__47___inst.ffx.TYPE = "#FF";
  defparam iSlice__47___inst.ffy.TYPE = "#FF";
  defparam iSlice__47___inst.fxmux.CONF = "F";
  defparam iSlice__47___inst.g.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__47___inst.gymux.CONF = "G";
  defparam iSlice__47___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__47___inst.ffy.INIT_VALUE = "LOW";
  defparam iSlice__47___inst.srffmux.CONF = "0";
  defparam iSlice__47___inst.srmux.CONF = "SR_B";
  defparam iSlice__47___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__47___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__47___inst.f.INIT = 16'h5;
  defparam iSlice__47___inst.g.INIT = 16'h5;
  SLICE iSlice__47___inst (
    .CIN(),
    .SR(net_rst_nInvLut_S1_SR_B_to_SR7_5_0),
    .CLK(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK7_5_0 ),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[0]_S1_F_B1_to_F17_5_0 ),
    .F2(net_U113_S1_F_B2_to_F27_5_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_Lut-U149_0_S1_G_B1_to_G17_5_0 ),
    .G2(net_U113_S1_G_B2_to_G27_5_0),
    .G3(),
    .G4(),
    .XQ(\net_cnt_lcd_reg[0]_XQ_to_S1_XQ7_5_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(\net_cnt_lcd_reg[1]_YQ_to_S1_YQ7_5_0 ),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__48___inst.f.CONF = "#LUT:D=((A3*~A2)*A1)";
  defparam iSlice__48___inst.fxmux.CONF = "F";
  defparam iSlice__48___inst.g.CONF = "#LUT:D=((A3*A2)*~A1)";
  defparam iSlice__48___inst.gymux.CONF = "G";
  defparam iSlice__48___inst.xused.CONF = "0";
  defparam iSlice__48___inst.yused.CONF = "0";
  defparam iSlice__48___inst.f.INIT = 16'h20;
  defparam iSlice__48___inst.g.INIT = 16'h40;
  SLICE iSlice__48___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_Lut-U224_0_0_S0_F_B1_to_F19_10_0 ),
    .F2(\net_cnt_lcd_reg[5]_S0_F_B2_to_F29_10_0 ),
    .F3(\net_cnt_lcd_reg[3]_S0_F_B3_to_F39_10_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[2]_S0_G_B1_to_G19_10_0 ),
    .G2(\net_cnt_lcd_reg[5]_S0_G_B2_to_G29_10_0 ),
    .G3(\net_cnt_lcd_reg[3]_S0_G_B3_to_G39_10_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U224_0_1_X_to_S0_X9_10_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U219_0_1_Y_to_S0_Y9_10_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__49___inst.f.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*A2)*~A1)+(((A4*A3)*~A2)*A1)+(((A4*A3)*~A2)*~A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*~A2)*A1)+(((~A4*~A3)*A2)*A1)";
  defparam iSlice__49___inst.fxmux.CONF = "F";
  defparam iSlice__49___inst.g.CONF = "#LUT:D=(((A4*A3)*A2)*A1)+(((A4*A3)*~A2)*A1)+(((A4*~A3)*A2)*A1)+(((A4*~A3)*A2)*~A1)+(((A4*~A3)*~A2)*A1)+(((A4*~A3)*~A2)*~A1)+(((~A4*A3)*A2)*A1)+(((~A4*A3)*A2)*~A1)+(((~A4*A3)*~A2)*A1)+(((~A4*~A3)*A2)*A1)+(((~A4*~A3)*A2)*~A1)+(((~A4*~A3)*~A2)*A1)+(((~A4*~A3)*~A2)*~A1)";
  defparam iSlice__49___inst.gymux.CONF = "G";
  defparam iSlice__49___inst.xused.CONF = "0";
  defparam iSlice__49___inst.yused.CONF = "0";
  defparam iSlice__49___inst.f.INIT = 16'hfda8;
  defparam iSlice__49___inst.g.INIT = 16'hafef;
  SLICE iSlice__49___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[1]_S0_F_B1_to_F17_10_0 ),
    .F2(\net_cnt_lcd_reg[3]_S0_F_B2_to_F27_10_0 ),
    .F3(\net_cnt_lcd_reg[5]_S0_F_B3_to_F37_10_0 ),
    .F4(\net_cnt_lcd_reg[2]_S0_F_B4_to_F47_10_0 ),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[2]_S0_G_B1_to_G17_10_0 ),
    .G2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G27_10_0 ),
    .G3(\net_cnt_lcd_reg[3]_S0_G_B3_to_G37_10_0 ),
    .G4(\net_cnt_lcd_reg[5]_S0_G_B4_to_G47_10_0 ),
    .XQ(),
    .X(\net_Lut-U129_0_X_to_S0_X7_10_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U154_0_Y_to_S0_Y7_10_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__50___inst.f.CONF = "#LUT:D=(((~A4*A3)*A2)*~A1)";
  defparam iSlice__50___inst.fxmux.CONF = "F";
  defparam iSlice__50___inst.g.CONF = "#LUT:D=1";
  defparam iSlice__50___inst.gymux.CONF = "G";
  defparam iSlice__50___inst.xused.CONF = "0";
  defparam iSlice__50___inst.yused.CONF = "0";
  defparam iSlice__50___inst.f.INIT = 16'h40;
  defparam iSlice__50___inst.g.INIT = 16'hffff;
  SLICE iSlice__50___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[2]_S1_F_B1_to_F111_10_0 ),
    .F2(\net_cnt_lcd_reg[5]_S1_F_B2_to_F211_10_0 ),
    .F3(\net_cnt_lcd_reg[3]_S1_F_B3_to_F311_10_0 ),
    .F4(\net_cnt_lcd_reg[1]_S1_F_B4_to_F411_10_0 ),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(\net_Lut-U216_0_0_X_to_S1_X11_10_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(net_U113_Y_to_S1_Y11_10_0),
    .YB(),
    .COUT()
  );

  defparam iSlice__51___inst.ckinv.CONF = "1";
  defparam iSlice__51___inst.dxmux.CONF = "1";
  defparam iSlice__51___inst.f.CONF = "#LUT:D=(A2*~A1)+(~A2*~A1)";
  defparam iSlice__51___inst.ffx.TYPE = "#FF";
  defparam iSlice__51___inst.fxmux.CONF = "F";
  defparam iSlice__51___inst.ffx.INIT_VALUE = "LOW";
  defparam iSlice__51___inst.srffmux.CONF = "0";
  defparam iSlice__51___inst.srmux.CONF = "SR_B";
  defparam iSlice__51___inst.ffx.SYNC_ATTR = "ASYNC";
  defparam iSlice__51___inst.ffy.SYNC_ATTR = "ASYNC";
  defparam iSlice__51___inst.f.INIT = 16'h5;
  SLICE iSlice__51___inst (
    .CIN(),
    .SR(net_rst_nInvLut_S1_SR_B_to_SR9_3_0),
    .CLK(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK9_3_0 ),
    .CE(),
    .BX(),
    .F1(\net_Lut-U115_1_S1_F_B1_to_F19_3_0 ),
    .F2(net_U113_S1_F_B2_to_F29_3_0),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(\net_lcd_db_reg[1]_XQ_to_S1_XQ9_3_0 ),
    .X(),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam iSlice__52___inst.f.CONF = "#LUT:D=(A2*~A1)";
  defparam iSlice__52___inst.fxmux.CONF = "F";
  defparam iSlice__52___inst.g.CONF = "#LUT:D=(A2*A1)+(~A2*~A1)";
  defparam iSlice__52___inst.gymux.CONF = "G";
  defparam iSlice__52___inst.xused.CONF = "0";
  defparam iSlice__52___inst.yused.CONF = "0";
  defparam iSlice__52___inst.f.INIT = 16'h4;
  defparam iSlice__52___inst.g.INIT = 16'h9;
  SLICE iSlice__52___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[6]_S0_F_B1_to_F17_5_0 ),
    .F2(\net_cnt_lcd_reg[0]_S0_F_B2_to_F27_5_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[0]_S0_G_B1_to_G17_5_0 ),
    .G2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G27_5_0 ),
    .G3(),
    .G4(),
    .XQ(),
    .X(\net_Lut-U232_0_0_X_to_S0_X7_5_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U149_0_Y_to_S0_Y7_5_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__53___inst.f.CONF = "#LUT:D=(~A2*~A1)";
  defparam iSlice__53___inst.fxmux.CONF = "F";
  defparam iSlice__53___inst.g.CONF = "#LUT:D=(A2*A1)";
  defparam iSlice__53___inst.gymux.CONF = "G";
  defparam iSlice__53___inst.xused.CONF = "0";
  defparam iSlice__53___inst.yused.CONF = "0";
  defparam iSlice__53___inst.f.INIT = 16'h1;
  defparam iSlice__53___inst.g.INIT = 16'h8;
  SLICE iSlice__53___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[1]_S1_F_B1_to_F111_9_0 ),
    .F2(\net_cnt_lcd_reg[2]_S1_F_B2_to_F211_9_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G111_9_0 ),
    .G2(\net_cnt_lcd_reg[5]_S1_G_B2_to_G211_9_0 ),
    .G3(),
    .G4(),
    .XQ(),
    .X(\net_Lut-U215_0_0_X_to_S1_X11_9_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U202_0_0_Y_to_S1_Y11_9_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__54___inst.f.CONF = "#LUT:D=(~A2*~A1)";
  defparam iSlice__54___inst.fxmux.CONF = "F";
  defparam iSlice__54___inst.g.CONF = "#LUT:D=(A2*A1)";
  defparam iSlice__54___inst.gymux.CONF = "G";
  defparam iSlice__54___inst.xused.CONF = "0";
  defparam iSlice__54___inst.yused.CONF = "0";
  defparam iSlice__54___inst.f.INIT = 16'h1;
  defparam iSlice__54___inst.g.INIT = 16'h8;
  SLICE iSlice__54___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[1]_S1_F_B1_to_F18_10_0 ),
    .F2(\net_cnt_lcd_reg[5]_S1_F_B2_to_F28_10_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[3]_S1_G_B1_to_G18_10_0 ),
    .G2(\net_cnt_lcd_reg[1]_S1_G_B2_to_G28_10_0 ),
    .G3(),
    .G4(),
    .XQ(),
    .X(\net_Lut-U177_0_0_X_to_S1_X8_10_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U226_0_0_Y_to_S1_Y8_10_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__55___inst.f.CONF = "#LUT:D=((~A3*A2)*A1)";
  defparam iSlice__55___inst.fxmux.CONF = "F";
  defparam iSlice__55___inst.g.CONF = "#LUT:D=((A3*A2)*A1)";
  defparam iSlice__55___inst.gymux.CONF = "G";
  defparam iSlice__55___inst.xused.CONF = "0";
  defparam iSlice__55___inst.yused.CONF = "0";
  defparam iSlice__55___inst.f.INIT = 16'h8;
  defparam iSlice__55___inst.g.INIT = 16'h80;
  SLICE iSlice__55___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[1]_S0_F_B1_to_F18_10_0 ),
    .F2(\net_cnt_lcd_reg[5]_S0_F_B2_to_F28_10_0 ),
    .F3(\net_cnt_lcd_reg[3]_S0_F_B3_to_F38_10_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S0_G_B1_to_G18_10_0 ),
    .G2(\net_cnt_lcd_reg[5]_S0_G_B2_to_G28_10_0 ),
    .G3(\net_cnt_lcd_reg[3]_S0_G_B3_to_G38_10_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U188_0_0_X_to_S0_X8_10_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U183_0_0_Y_to_S0_Y8_10_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__56___inst.f.CONF = "#LUT:D=(A2*~A1)";
  defparam iSlice__56___inst.fxmux.CONF = "F";
  defparam iSlice__56___inst.g.CONF = "#LUT:D=(A2*~A1)";
  defparam iSlice__56___inst.gymux.CONF = "G";
  defparam iSlice__56___inst.xused.CONF = "0";
  defparam iSlice__56___inst.yused.CONF = "0";
  defparam iSlice__56___inst.f.INIT = 16'h4;
  defparam iSlice__56___inst.g.INIT = 16'h4;
  SLICE iSlice__56___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[5]_S1_F_B1_to_F110_9_0 ),
    .F2(\net_cnt_lcd_reg[3]_S1_F_B2_to_F210_9_0 ),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G110_9_0 ),
    .G2(\net_cnt_lcd_reg[3]_S1_G_B2_to_G210_9_0 ),
    .G3(),
    .G4(),
    .XQ(),
    .X(\net_Lut-U227_0_X_to_S1_X10_9_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U161_0_0_Y_to_S1_Y10_9_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__57___inst.f.CONF = "#LUT:D=((A3*~A2)*~A1)";
  defparam iSlice__57___inst.fxmux.CONF = "F";
  defparam iSlice__57___inst.g.CONF = "#LUT:D=((A3*~A2)*~A1)";
  defparam iSlice__57___inst.gymux.CONF = "G";
  defparam iSlice__57___inst.xused.CONF = "0";
  defparam iSlice__57___inst.yused.CONF = "0";
  defparam iSlice__57___inst.f.INIT = 16'h10;
  defparam iSlice__57___inst.g.INIT = 16'h10;
  SLICE iSlice__57___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(\net_cnt_lcd_reg[1]_S1_F_B1_to_F18_6_0 ),
    .F2(\net_cnt_lcd_reg[3]_S1_F_B2_to_F28_6_0 ),
    .F3(\net_cnt_lcd_reg[5]_S1_F_B3_to_F38_6_0 ),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G18_6_0 ),
    .G2(\net_cnt_lcd_reg[5]_S1_G_B2_to_G28_6_0 ),
    .G3(\net_cnt_lcd_reg[3]_S1_G_B3_to_G38_6_0 ),
    .G4(),
    .XQ(),
    .X(\net_Lut-U190_0_1_X_to_S1_X8_6_0 ),
    .F5(),
    .XB(),
    .YQ(),
    .Y(\net_Lut-U186_0_Y_to_S1_Y8_6_0 ),
    .YB(),
    .COUT()
  );

  defparam iSlice__58___inst.f.CONF = "#LUT:D=0";
  defparam iSlice__58___inst.fxmux.CONF = "F";
  defparam iSlice__58___inst.xused.CONF = "0";
  defparam iSlice__58___inst.f.INIT = 16'h0;
  SLICE iSlice__58___inst (
    .CIN(),
    .SR(),
    .CLK(),
    .CE(),
    .BX(),
    .F1(),
    .F2(),
    .F3(),
    .F4(),
    .F5IN(),
    .BY(),
    .G1(),
    .G2(),
    .G3(),
    .G4(),
    .XQ(),
    .X(net_U108_X_to_S0_X6_3_0),
    .F5(),
    .XB(),
    .YQ(),
    .Y(),
    .YB(),
    .COUT()
  );

  defparam \lcd_db[6]_inst .driveattrbox.CONF = "12";
  defparam \lcd_db[6]_inst .ioattrbox.CONF = "LVTTL";
  defparam \lcd_db[6]_inst .omux.CONF = "O";
  defparam \lcd_db[6]_inst .outmux.CONF = "1";
  defparam \lcd_db[6]_inst .slew.CONF = "SLOW";
  IOB \lcd_db[6]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_lcd_db_reg[6]_LEFT_O2_to_OUT9_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_db[6])
  );

  defparam \lcd_db[5]_inst .driveattrbox.CONF = "12";
  defparam \lcd_db[5]_inst .ioattrbox.CONF = "LVTTL";
  defparam \lcd_db[5]_inst .omux.CONF = "O";
  defparam \lcd_db[5]_inst .outmux.CONF = "1";
  defparam \lcd_db[5]_inst .slew.CONF = "SLOW";
  IOB \lcd_db[5]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_lcd_db_reg[5]_LEFT_O3_to_OUT9_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_db[5])
  );

  defparam \lcd_db[4]_inst .driveattrbox.CONF = "12";
  defparam \lcd_db[4]_inst .ioattrbox.CONF = "LVTTL";
  defparam \lcd_db[4]_inst .omux.CONF = "O";
  defparam \lcd_db[4]_inst .outmux.CONF = "1";
  defparam \lcd_db[4]_inst .slew.CONF = "SLOW";
  IOB \lcd_db[4]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_lcd_db_reg[4]_LEFT_O1_to_OUT10_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_db[4])
  );

  defparam \lcd_db[3]_inst .driveattrbox.CONF = "12";
  defparam \lcd_db[3]_inst .ioattrbox.CONF = "LVTTL";
  defparam \lcd_db[3]_inst .omux.CONF = "O";
  defparam \lcd_db[3]_inst .outmux.CONF = "1";
  defparam \lcd_db[3]_inst .slew.CONF = "SLOW";
  IOB \lcd_db[3]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_lcd_db_reg[3]_LEFT_O2_to_OUT10_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_db[3])
  );

  defparam \lcd_db[2]_inst .driveattrbox.CONF = "12";
  defparam \lcd_db[2]_inst .ioattrbox.CONF = "LVTTL";
  defparam \lcd_db[2]_inst .omux.CONF = "O";
  defparam \lcd_db[2]_inst .outmux.CONF = "1";
  defparam \lcd_db[2]_inst .slew.CONF = "SLOW";
  IOB \lcd_db[2]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_lcd_db_reg[2]_LEFT_O1_to_OUT8_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_db[2])
  );

  defparam \lcd_db[1]_inst .driveattrbox.CONF = "12";
  defparam \lcd_db[1]_inst .ioattrbox.CONF = "LVTTL";
  defparam \lcd_db[1]_inst .omux.CONF = "O";
  defparam \lcd_db[1]_inst .outmux.CONF = "1";
  defparam \lcd_db[1]_inst .slew.CONF = "SLOW";
  IOB \lcd_db[1]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_lcd_db_reg[1]_LEFT_O1_to_OUT9_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_db[1])
  );

  defparam \lcd_db[0]_inst .driveattrbox.CONF = "12";
  defparam \lcd_db[0]_inst .ioattrbox.CONF = "LVTTL";
  defparam \lcd_db[0]_inst .omux.CONF = "O";
  defparam \lcd_db[0]_inst .outmux.CONF = "1";
  defparam \lcd_db[0]_inst .slew.CONF = "SLOW";
  IOB \lcd_db[0]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(\net_lcd_db_reg[0]_LEFT_O1_to_OUT4_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_db[0])
  );

  defparam rst_n_inst.imux.CONF = "1";
  defparam rst_n_inst.ioattrbox.CONF = "LVTTL";
  IOB rst_n_inst (
    .TRI(),
    .TRICE(),
    .OUT(),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(\net_Buf-pad-rst_n_IN_to_RIGHT_I35_54_0 ),
    .IQ(),
    .PAD(rst_n)
  );

  defparam \lcd_db[7]_inst .driveattrbox.CONF = "12";
  defparam \lcd_db[7]_inst .ioattrbox.CONF = "LVTTL";
  defparam \lcd_db[7]_inst .omux.CONF = "O";
  defparam \lcd_db[7]_inst .outmux.CONF = "1";
  defparam \lcd_db[7]_inst .slew.CONF = "SLOW";
  IOB \lcd_db[7]_inst  (
    .TRI(),
    .TRICE(),
    .OUT(net_U108_LEFT_O1_to_OUT14_2_0),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_db[7])
  );

  defparam lcd_rw_inst.driveattrbox.CONF = "12";
  defparam lcd_rw_inst.ioattrbox.CONF = "LVTTL";
  defparam lcd_rw_inst.omux.CONF = "O";
  defparam lcd_rw_inst.outmux.CONF = "1";
  defparam lcd_rw_inst.slew.CONF = "SLOW";
  IOB lcd_rw_inst (
    .TRI(),
    .TRICE(),
    .OUT(net_U108_LEFT_O3_to_OUT5_2_0),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_rw)
  );

  defparam lcd_rst_inst.driveattrbox.CONF = "12";
  defparam lcd_rst_inst.ioattrbox.CONF = "LVTTL";
  defparam lcd_rst_inst.omux.CONF = "O";
  defparam lcd_rst_inst.outmux.CONF = "1";
  defparam lcd_rst_inst.slew.CONF = "SLOW";
  IOB lcd_rst_inst (
    .TRI(),
    .TRICE(),
    .OUT(\net_Buf-pad-rst_n_LEFT_O3_to_OUT13_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_rst)
  );

  defparam lcd_en_inst.driveattrbox.CONF = "12";
  defparam lcd_en_inst.ioattrbox.CONF = "LVTTL";
  defparam lcd_en_inst.omux.CONF = "O";
  defparam lcd_en_inst.outmux.CONF = "1";
  defparam lcd_en_inst.slew.CONF = "SLOW";
  IOB lcd_en_inst (
    .TRI(),
    .TRICE(),
    .OUT(\net_Lut-U232_0_0_LEFT_O2_to_OUT6_2_0 ),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_en)
  );

  defparam lcd_rs_inst.driveattrbox.CONF = "12";
  defparam lcd_rs_inst.ioattrbox.CONF = "LVTTL";
  defparam lcd_rs_inst.omux.CONF = "O";
  defparam lcd_rs_inst.outmux.CONF = "1";
  defparam lcd_rs_inst.slew.CONF = "SLOW";
  IOB lcd_rs_inst (
    .TRI(),
    .TRICE(),
    .OUT(net_U113_LEFT_O1_to_OUT6_2_0),
    .OUTCE(),
    .INCE(),
    .CLK(),
    .SR(),
    .IN(),
    .IQ(),
    .PAD(lcd_rs)
  );

  defparam iGclk_buf__0___inst.cemux.CONF = "1";
  defparam iGclk_buf__0___inst.disable_attr.CONF = "LOW";
  GCLK iGclk_buf__0___inst (
    .CE(),
    .IN(\net_Buf-pad-clk_CLKB_GCLKBUF1_IN_to_IN35_28_0 ),
    .OUT(\net_IBuf-clkpad-clk_OUT_to_CLKB_GCLK1_PW35_28_0 )
  );

  defparam clk_inst.ioattrbox.CONF = "LVTTL";
  GCLKIOB clk_inst (
    .PAD(clk),
    .GCLKOUT(\net_Buf-pad-clk_GCLKOUT_to_CLKB_CLKPAD135_28_0 )
  );

  defparam GSB_CNT_7_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e14.CONF = "0";
  defparam GSB_CNT_7_6_0_inst.sps_e15.CONF = "01";
  defparam GSB_CNT_7_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_e17.CONF = "10";
  defparam GSB_CNT_7_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_e2.CONF = "0";
  defparam GSB_CNT_7_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e3.CONF = "10";
  defparam GSB_CNT_7_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_e8.CONF = "0";
  defparam GSB_CNT_7_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_h6e0.CONF = "0001";
  defparam GSB_CNT_7_6_0_inst.sps_h6e1.CONF = "0001";
  defparam GSB_CNT_7_6_0_inst.sps_h6e11.CONF = "001";
  defparam GSB_CNT_7_6_0_inst.sps_h6e2.CONF = "0001";
  defparam GSB_CNT_7_6_0_inst.sps_h6e3.CONF = "0001";
  defparam GSB_CNT_7_6_0_inst.sps_h6e5.CONF = "001";
  defparam GSB_CNT_7_6_0_inst.sps_h6e7.CONF = "001";
  defparam GSB_CNT_7_6_0_inst.sps_h6e9.CONF = "001";
  defparam GSB_CNT_7_6_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_6_0_inst.sps_h6w1.CONF = "0010";
  defparam GSB_CNT_7_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_6_0_inst.sps_h6w2.CONF = "0010";
  defparam GSB_CNT_7_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_6_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_llh6.CONF = "00";
  defparam GSB_CNT_7_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_6_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_out0.CONF = "001110";
  defparam GSB_CNT_7_6_0_inst.sps_out1.CONF = "001110";
  defparam GSB_CNT_7_6_0_inst.sps_out2.CONF = "001101";
  defparam GSB_CNT_7_6_0_inst.sps_out3.CONF = "001101";
  defparam GSB_CNT_7_6_0_inst.sps_out4.CONF = "100111";
  defparam GSB_CNT_7_6_0_inst.sps_out5.CONF = "101011";
  defparam GSB_CNT_7_6_0_inst.sps_out6.CONF = "001110";
  defparam GSB_CNT_7_6_0_inst.sps_out7.CONF = "101011";
  defparam GSB_CNT_7_6_0_inst.sps_s0.CONF = "0";
  defparam GSB_CNT_7_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_7_6_0_inst.sps_s0_f_b1.CONF = "011111011";
  defparam GSB_CNT_7_6_0_inst.sps_s0_f_b2.CONF = "001111110";
  defparam GSB_CNT_7_6_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_6_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_6_0_inst.sps_s0_g_b1.CONF = "100101";
  defparam GSB_CNT_7_6_0_inst.sps_s0_g_b2.CONF = "001000";
  defparam GSB_CNT_7_6_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_s0_sr_b.CONF = "011011";
  defparam GSB_CNT_7_6_0_inst.sps_s1.CONF = "10";
  defparam GSB_CNT_7_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_s12.CONF = "0";
  defparam GSB_CNT_7_6_0_inst.sps_s13.CONF = "10";
  defparam GSB_CNT_7_6_0_inst.sps_s14.CONF = "01";
  defparam GSB_CNT_7_6_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_s17.CONF = "10";
  defparam GSB_CNT_7_6_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_s1_clk_b.CONF = "101011";
  defparam GSB_CNT_7_6_0_inst.sps_s1_f_b1.CONF = "001111101";
  defparam GSB_CNT_7_6_0_inst.sps_s1_f_b2.CONF = "011111011";
  defparam GSB_CNT_7_6_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_6_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_6_0_inst.sps_s1_g_b1.CONF = "011000";
  defparam GSB_CNT_7_6_0_inst.sps_s1_g_b2.CONF = "011101";
  defparam GSB_CNT_7_6_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_s1_sr_b.CONF = "011011";
  defparam GSB_CNT_7_6_0_inst.sps_s2.CONF = "01";
  defparam GSB_CNT_7_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_s5.CONF = "10";
  defparam GSB_CNT_7_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_s7.CONF = "0";
  defparam GSB_CNT_7_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_6_0_inst.sps_v6n0.CONF = "0001";
  defparam GSB_CNT_7_6_0_inst.sps_v6n1.CONF = "0001";
  defparam GSB_CNT_7_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_6_0_inst.sps_v6n2.CONF = "0011";
  defparam GSB_CNT_7_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_6_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_6_0_inst.sps_v6s0.CONF = "0000";
  defparam GSB_CNT_7_6_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_7_6_0_inst.sps_v6s10.CONF = "001";
  defparam GSB_CNT_7_6_0_inst.sps_v6s2.CONF = "0000";
  defparam GSB_CNT_7_6_0_inst.sps_v6s3.CONF = "0000";
  defparam GSB_CNT_7_6_0_inst.sps_v6s4.CONF = "001";
  defparam GSB_CNT_7_6_0_inst.sps_v6s6.CONF = "001";
  defparam GSB_CNT_7_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w19.CONF = "0";
  defparam GSB_CNT_7_6_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e5_w5.CONF = "0";
  defparam GSB_CNT_7_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n14_e10.CONF = "0";
  defparam GSB_CNT_7_6_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s3_w5.CONF = "0";
  defparam GSB_CNT_7_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_6_0_inst (
    .E0(),
    .E1(),
    .E2(\net_cnt_lcd_reg[5]_E2_to_W27_7_0 ),
    .E3(\net_cnt_lcd_reg[5]_E3_to_W37_7_0 ),
    .E4(),
    .E5(\net_cnt_lcd_reg[1]_E5_to_W57_7_0 ),
    .E6(),
    .E7(),
    .E8(\net_cnt_lcd_reg[4]_E8_to_W87_7_0 ),
    .E9(),
    .E10(\net_Lut-U141_0_W10_to_E107_6_0 ),
    .E11(),
    .E12(),
    .E13(),
    .E14(\net_cnt_lcd_reg[6]_E14_to_W147_7_0 ),
    .E15(\net_cnt_lcd_reg[7]_E15_to_W157_7_0 ),
    .E16(),
    .E17(\net_cnt_lcd_reg[7]_E17_to_W177_7_0 ),
    .E18(),
    .E19(\net_Lut-U138_0_W19_to_E197_6_0 ),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(net_rst_nInvLut_S8_to_N87_6_0),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(\net_cnt_lcd_reg[1]_E5_to_W57_6_0 ),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(\net_cnt_lcd_reg[6]_W19_to_E197_5_0 ),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(\net_cnt_lcd_reg[5]_S0_to_N08_6_0 ),
    .S1(\net_cnt_lcd_reg[5]_S1_to_N18_6_0 ),
    .S2(\net_cnt_lcd_reg[5]_S2_to_N28_6_0 ),
    .S3(\net_cnt_lcd_reg[1]_S3_to_N38_6_0 ),
    .S4(net_U113_N4_to_S47_6_0),
    .S5(\net_cnt_lcd_reg[4]_S5_to_N58_6_0 ),
    .S6(\net_Lut-U143_0_N6_to_S67_6_0 ),
    .S7(\net_cnt_lcd_reg[4]_S7_to_N78_6_0 ),
    .S8(),
    .S9(\net_Lut-U136_0_N9_to_S97_6_0 ),
    .S10(),
    .S11(),
    .S12(\net_cnt_lcd_reg[7]_S12_to_N128_6_0 ),
    .S13(\net_cnt_lcd_reg[6]_S13_to_N138_6_0 ),
    .S14(\net_cnt_lcd_reg[7]_S14_to_N148_6_0 ),
    .S15(net_U113_N15_to_S157_6_0),
    .S16(),
    .S17(\net_cnt_lcd_reg[5]_S17_to_N178_6_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(\net_cnt_lcd_reg[5]_H6E0_to_H6M07_9_0 ),
    .H6E1(\net_cnt_lcd_reg[4]_H6E1_to_H6W17_12_0 ),
    .H6E2(\net_cnt_lcd_reg[7]_H6E2_to_H6M27_9_0 ),
    .H6E3(\net_cnt_lcd_reg[6]_H6E3_to_H6M37_9_0 ),
    .H6E4(),
    .H6E5(\net_cnt_lcd_reg[5]_H6E5_to_H6M57_9_0 ),
    .H6E6(),
    .H6E7(\net_cnt_lcd_reg[6]_H6E7_to_H6M77_9_0 ),
    .H6E8(),
    .H6E9(\net_cnt_lcd_reg[4]_H6E9_to_H6W97_12_0 ),
    .H6E10(),
    .H6E11(\net_cnt_lcd_reg[5]_H6E11_to_H6M117_9_0 ),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_cnt_lcd_reg[4]_H6W1_to_H6M17_3_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBB1_to_GCLK17_3_0 ),
    .GCLK0(),
    .OUT0(\net_cnt_lcd_reg[5]_OUT0_to_OUT_W07_7_0 ),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(\net_cnt_lcd_reg[4]_V6N1_to_V6M14_6_0 ),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(\net_cnt_lcd_reg[5]_V6S0_to_V6M010_6_0 ),
    .V6S1(),
    .V6S2(\net_cnt_lcd_reg[6]_V6S2_to_V6M210_6_0 ),
    .V6S3(\net_cnt_lcd_reg[5]_V6S3_to_V6M310_6_0 ),
    .V6S4(\net_cnt_lcd_reg[5]_V6S4_to_V6M410_6_0 ),
    .V6S5(),
    .V6S6(\net_cnt_lcd_reg[7]_V6S6_to_V6M610_6_0 ),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(\net_cnt_lcd_reg[7]_V6S10_to_V6M1010_6_0 ),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U143_0_S0_F_B1_to_F17_6_0 ),
    .S0_F_B2(net_U113_S0_F_B2_to_F27_6_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Lut-U141_0_S0_G_B1_to_G17_6_0 ),
    .S0_G_B2(net_U113_S0_G_B2_to_G27_6_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK7_6_0 ),
    .S0_SR_B(net_rst_nInvLut_S0_SR_B_to_SR7_6_0),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_cnt_lcd_reg[4]_XQ_to_S0_XQ7_6_0 ),
    .S0_YQ(\net_cnt_lcd_reg[5]_YQ_to_S0_YQ7_6_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U138_0_S1_F_B1_to_F17_6_0 ),
    .S1_F_B2(net_U113_S1_F_B2_to_F27_6_0),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(\net_Lut-U136_0_S1_G_B1_to_G17_6_0 ),
    .S1_G_B2(net_U113_S1_G_B2_to_G27_6_0),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK7_6_0 ),
    .S1_SR_B(net_rst_nInvLut_S1_SR_B_to_SR7_6_0),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(\net_cnt_lcd_reg[6]_XQ_to_S1_XQ7_6_0 ),
    .S1_YQ(\net_cnt_lcd_reg[7]_YQ_to_S1_YQ7_6_0 ),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_9_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_e21.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_e9.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_9_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_9_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n10.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_n16.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.sps_n17.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n23.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_n4.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_out0.CONF = "000111";
  defparam GSB_CNT_7_9_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_out2.CONF = "000111";
  defparam GSB_CNT_7_9_0_inst.sps_out3.CONF = "000111";
  defparam GSB_CNT_7_9_0_inst.sps_out4.CONF = "000111";
  defparam GSB_CNT_7_9_0_inst.sps_out5.CONF = "001011";
  defparam GSB_CNT_7_9_0_inst.sps_out6.CONF = "011110";
  defparam GSB_CNT_7_9_0_inst.sps_out7.CONF = "011101";
  defparam GSB_CNT_7_9_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_s0_f_b1.CONF = "100011111";
  defparam GSB_CNT_7_9_0_inst.sps_s0_f_b2.CONF = "010101111";
  defparam GSB_CNT_7_9_0_inst.sps_s0_f_b3.CONF = "100111101";
  defparam GSB_CNT_7_9_0_inst.sps_s0_f_b4.CONF = "011011111";
  defparam GSB_CNT_7_9_0_inst.sps_s0_g_b1.CONF = "100100";
  defparam GSB_CNT_7_9_0_inst.sps_s0_g_b2.CONF = "010011";
  defparam GSB_CNT_7_9_0_inst.sps_s0_g_b3.CONF = "010000";
  defparam GSB_CNT_7_9_0_inst.sps_s0_g_b4.CONF = "010011";
  defparam GSB_CNT_7_9_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s18.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_s1_f_b1.CONF = "001110111";
  defparam GSB_CNT_7_9_0_inst.sps_s1_f_b2.CONF = "100111110";
  defparam GSB_CNT_7_9_0_inst.sps_s1_f_b3.CONF = "011011111";
  defparam GSB_CNT_7_9_0_inst.sps_s1_f_b4.CONF = "011110111";
  defparam GSB_CNT_7_9_0_inst.sps_s1_g_b1.CONF = "110111";
  defparam GSB_CNT_7_9_0_inst.sps_s1_g_b2.CONF = "001111";
  defparam GSB_CNT_7_9_0_inst.sps_s1_g_b3.CONF = "010010";
  defparam GSB_CNT_7_9_0_inst.sps_s1_g_b4.CONF = "010010";
  defparam GSB_CNT_7_9_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s4.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s6.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_s9.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_9_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_v6n1.CONF = "0100";
  defparam GSB_CNT_7_9_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_v6n3.CONF = "0100";
  defparam GSB_CNT_7_9_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_9_0_inst.sps_v6s0.CONF = "0000";
  defparam GSB_CNT_7_9_0_inst.sps_v6s1.CONF = "0000";
  defparam GSB_CNT_7_9_0_inst.sps_v6s10.CONF = "011";
  defparam GSB_CNT_7_9_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_9_0_inst.sps_v6s4.CONF = "011";
  defparam GSB_CNT_7_9_0_inst.sps_v6s6.CONF = "011";
  defparam GSB_CNT_7_9_0_inst.sps_v6s8.CONF = "001";
  defparam GSB_CNT_7_9_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w16.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w19.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w23.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_9_0_inst.sps_w9.CONF = "10";
  defparam GSB_CNT_7_9_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n10_e6.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n16_e12.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n17_e17.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n19_e19.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n1_w2.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n23_e23.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s17_n17.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s1_w7.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s4_e2.CONF = "0";
  defparam GSB_CNT_7_9_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_9_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_9_0_inst (
    .E0(),
    .E1(),
    .E2(\net_cnt_lcd_reg[5]_E2_to_W27_10_0 ),
    .E3(),
    .E4(),
    .E5(),
    .E6(\net_cnt_lcd_reg[4]_E6_to_W67_10_0 ),
    .E7(),
    .E8(),
    .E9(\net_cnt_lcd_reg[4]_E9_to_W97_10_0 ),
    .E10(),
    .E11(),
    .E12(\net_cnt_lcd_reg[7]_E12_to_W127_10_0 ),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(\net_cnt_lcd_reg[6]_E17_to_W177_10_0 ),
    .E18(),
    .E19(\net_Lut-U229_0_W19_to_E197_9_0 ),
    .E20(),
    .E21(),
    .E22(),
    .E23(\net_cnt_lcd_reg[5]_E23_to_W237_10_0 ),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(\net_cnt_lcd_reg[2]_S20_to_N207_9_0 ),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(\net_cnt_lcd_reg[0]_E2_to_W27_9_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(\net_Lut-U176_0_1_W7_to_E77_8_0 ),
    .W8(),
    .W9(\net_Lut-U201_0_0_W9_to_E97_8_0 ),
    .W10(),
    .W11(\net_Lut-U189_2_E11_to_W117_9_0 ),
    .W12(),
    .W13(),
    .W14(\net_cnt_lcd_reg[3]_E14_to_W147_9_0 ),
    .W15(\net_cnt_lcd_reg[7]_E15_to_W157_9_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(\net_Lut-U201_0_0_W19_to_E197_8_0 ),
    .W20(\net_cnt_lcd_reg[1]_E20_to_W207_9_0 ),
    .W21(\net_cnt_lcd_reg[0]_E21_to_W217_9_0 ),
    .W22(),
    .W23(\net_Lut-U130_0_1_W23_to_E237_8_0 ),
    .S0(\net_Lut-U176_0_1_N0_to_S07_9_0 ),
    .S1(\net_Lut-U176_0_1_N1_to_S17_9_0 ),
    .S2(),
    .S3(),
    .S4(\net_cnt_lcd_reg[5]_S4_to_N48_9_0 ),
    .S5(),
    .S6(\net_cnt_lcd_reg[5]_S6_to_N68_9_0 ),
    .S7(),
    .S8(),
    .S9(\net_cnt_lcd_reg[4]_S9_to_N98_9_0 ),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(\net_cnt_lcd_reg[6]_S17_to_N178_9_0 ),
    .S18(\net_cnt_lcd_reg[7]_S18_to_N188_9_0 ),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(\net_cnt_lcd_reg[5]_H6E0_to_H6M07_9_0 ),
    .H6M1(\net_cnt_lcd_reg[4]_H6E1_to_H6W17_12_0 ),
    .H6M2(\net_cnt_lcd_reg[7]_H6E2_to_H6M27_9_0 ),
    .H6M3(\net_cnt_lcd_reg[6]_H6E3_to_H6M37_9_0 ),
    .H6M4(),
    .H6M5(\net_cnt_lcd_reg[5]_H6E5_to_H6M57_9_0 ),
    .H6M6(),
    .H6M7(\net_cnt_lcd_reg[6]_H6E7_to_H6M77_9_0 ),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(\net_cnt_lcd_reg[5]_H6E11_to_H6M117_9_0 ),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(\net_Lut-U127_0_OUT6_to_OUT_E67_8_0 ),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(\net_Lut-U127_0_0_OUT6_to_OUT_E67_9_0 ),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(\net_Lut-U201_0_0_V6S0_to_V6M010_9_0 ),
    .V6S1(\net_Lut-U201_0_0_V6S1_to_V6M110_9_0 ),
    .V6S2(),
    .V6S3(),
    .V6S4(\net_cnt_lcd_reg[5]_V6S4_to_V6M410_9_0 ),
    .V6S5(),
    .V6S6(\net_cnt_lcd_reg[6]_V6S6_to_V6M610_9_0 ),
    .V6S7(),
    .V6S8(\net_Lut-U201_0_0_V6S8_to_V6M810_9_0 ),
    .V6S9(),
    .V6S10(\net_cnt_lcd_reg[5]_V6S10_to_V6M1010_9_0 ),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[2]_S0_F_B1_to_F17_9_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[7]_S0_F_B2_to_F27_9_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[6]_S0_F_B3_to_F37_9_0 ),
    .S0_F_B4(\net_cnt_lcd_reg[0]_S0_F_B4_to_F47_9_0 ),
    .S0_G_B1(\net_cnt_lcd_reg[2]_S0_G_B1_to_G17_9_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G27_9_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[5]_S0_G_B3_to_G37_9_0 ),
    .S0_G_B4(\net_cnt_lcd_reg[3]_S0_G_B4_to_G47_9_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U201_0_0_X_to_S0_X7_9_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U132_0_Y_to_S0_Y7_9_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U189_2_S1_F_B1_to_F17_9_0 ),
    .S1_F_B2(\net_Lut-U176_0_1_S1_F_B2_to_F27_9_0 ),
    .S1_F_B3(\net_Lut-U132_0_S1_F_B3_to_F37_9_0 ),
    .S1_F_B4(\net_Lut-U229_0_S1_F_B4_to_F47_9_0 ),
    .S1_G_B1(\net_Lut-U127_0_0_S1_G_B1_to_G17_9_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[7]_S1_G_B2_to_G27_9_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[6]_S1_G_B3_to_G37_9_0 ),
    .S1_G_B4(\net_cnt_lcd_reg[0]_S1_G_B4_to_G47_9_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U130_0_1_X_to_S1_X7_9_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U127_0_Y_to_S1_Y7_9_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_7_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_h6w6.CONF = "000";
  defparam GSB_CNT_7_7_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_7_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_7_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_out0.CONF = "000111";
  defparam GSB_CNT_7_7_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_out2.CONF = "001011";
  defparam GSB_CNT_7_7_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_7_7_0_inst.sps_out4.CONF = "011110";
  defparam GSB_CNT_7_7_0_inst.sps_out5.CONF = "001011";
  defparam GSB_CNT_7_7_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s0_f_b1.CONF = "011111110";
  defparam GSB_CNT_7_7_0_inst.sps_s0_f_b2.CONF = "110111111";
  defparam GSB_CNT_7_7_0_inst.sps_s0_f_b3.CONF = "001110111";
  defparam GSB_CNT_7_7_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_7_0_inst.sps_s0_g_b1.CONF = "100000";
  defparam GSB_CNT_7_7_0_inst.sps_s0_g_b2.CONF = "100111";
  defparam GSB_CNT_7_7_0_inst.sps_s0_g_b3.CONF = "011100";
  defparam GSB_CNT_7_7_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s18.CONF = "10";
  defparam GSB_CNT_7_7_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s1_f_b1.CONF = "010011111";
  defparam GSB_CNT_7_7_0_inst.sps_s1_f_b2.CONF = "010101111";
  defparam GSB_CNT_7_7_0_inst.sps_s1_f_b3.CONF = "010111011";
  defparam GSB_CNT_7_7_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_7_0_inst.sps_s1_g_b1.CONF = "011000";
  defparam GSB_CNT_7_7_0_inst.sps_s1_g_b2.CONF = "100011";
  defparam GSB_CNT_7_7_0_inst.sps_s1_g_b3.CONF = "100011";
  defparam GSB_CNT_7_7_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s5.CONF = "10";
  defparam GSB_CNT_7_7_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_7_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_v6s1.CONF = "0000";
  defparam GSB_CNT_7_7_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_7_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_v6s6.CONF = "001";
  defparam GSB_CNT_7_7_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_7_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_w10.CONF = "10";
  defparam GSB_CNT_7_7_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_7_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e14_w14.CONF = "0";
  defparam GSB_CNT_7_7_0_inst.switch_e15_w15.CONF = "0";
  defparam GSB_CNT_7_7_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e19_w19.CONF = "0";
  defparam GSB_CNT_7_7_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e2_w2.CONF = "0";
  defparam GSB_CNT_7_7_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_e8_w8.CONF = "0";
  defparam GSB_CNT_7_7_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_n9_e9.CONF = "0";
  defparam GSB_CNT_7_7_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s10_w8.CONF = "0";
  defparam GSB_CNT_7_7_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s15_w17.CONF = "0";
  defparam GSB_CNT_7_7_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_7_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_7_0_inst (
    .E0(),
    .E1(),
    .E2(\net_cnt_lcd_reg[5]_E2_to_W27_8_0 ),
    .E3(\net_Lut-U178_0_W3_to_E37_7_0 ),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(\net_cnt_lcd_reg[4]_E8_to_W87_8_0 ),
    .E9(\net_Lut-U201_0_0_W9_to_E97_7_0 ),
    .E10(),
    .E11(\net_Lut-U174_0_W11_to_E117_7_0 ),
    .E12(),
    .E13(),
    .E14(\net_cnt_lcd_reg[6]_E14_to_W147_8_0 ),
    .E15(\net_cnt_lcd_reg[7]_E15_to_W157_8_0 ),
    .E16(),
    .E17(),
    .E18(),
    .E19(\net_Lut-U138_0_W19_to_E197_7_0 ),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(\net_cnt_lcd_reg[2]_S6_to_N67_7_0 ),
    .N7(),
    .N8(\net_Lut-U144_0_0_S8_to_N87_7_0 ),
    .N9(),
    .N10(),
    .N11(\net_cnt_lcd_reg[3]_S11_to_N117_7_0 ),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(\net_cnt_lcd_reg[3]_S18_to_N187_7_0 ),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(\net_cnt_lcd_reg[5]_E2_to_W27_7_0 ),
    .W3(\net_cnt_lcd_reg[5]_E3_to_W37_7_0 ),
    .W4(),
    .W5(\net_cnt_lcd_reg[1]_E5_to_W57_7_0 ),
    .W6(),
    .W7(),
    .W8(\net_cnt_lcd_reg[4]_E8_to_W87_7_0 ),
    .W9(),
    .W10(\net_Lut-U141_0_W10_to_E107_6_0 ),
    .W11(),
    .W12(),
    .W13(),
    .W14(\net_cnt_lcd_reg[6]_E14_to_W147_7_0 ),
    .W15(\net_cnt_lcd_reg[7]_E15_to_W157_7_0 ),
    .W16(),
    .W17(\net_cnt_lcd_reg[7]_E17_to_W177_7_0 ),
    .W18(),
    .W19(\net_Lut-U138_0_W19_to_E197_6_0 ),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(\net_Lut-U205_0_0_S5_to_N58_7_0 ),
    .S6(),
    .S7(),
    .S8(),
    .S9(\net_Lut-U191_1_N9_to_S97_7_0 ),
    .S10(\net_cnt_lcd_reg[4]_S10_to_N108_7_0 ),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(\net_cnt_lcd_reg[7]_S15_to_N158_7_0 ),
    .S16(),
    .S17(),
    .S18(\net_Lut-U225_0_S18_to_N188_7_0 ),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(\net_Lut-U225_0_H6W2_to_H6M27_7_0 ),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_Lut-U173_1_H6W6_to_H6M67_4_0 ),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(\net_Lut-U175_0_0_OUT0_to_OUT_W07_8_0 ),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(\net_cnt_lcd_reg[5]_OUT0_to_OUT_W07_7_0 ),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(\net_Lut-U205_0_0_V6S1_to_V6M110_7_0 ),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(\net_Lut-U205_0_0_V6S6_to_V6M610_7_0 ),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U201_0_0_S0_F_B1_to_F17_7_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[5]_S0_F_B2_to_F27_7_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[3]_S0_F_B3_to_F37_7_0 ),
    .S0_F_B4(),
    .S0_G_B1(\net_cnt_lcd_reg[1]_S0_G_B1_to_G17_7_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[3]_S0_G_B2_to_G27_7_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[2]_S0_G_B3_to_G37_7_0 ),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U175_0_0_X_to_S0_X7_7_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U205_0_0_Y_to_S0_Y7_7_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[5]_S1_F_B1_to_F17_7_0 ),
    .S1_F_B2(\net_Lut-U144_0_0_S1_F_B2_to_F27_7_0 ),
    .S1_F_B3(\net_cnt_lcd_reg[4]_S1_F_B3_to_F37_7_0 ),
    .S1_F_B4(),
    .S1_G_B1(\net_Lut-U191_1_S1_G_B1_to_G17_7_0 ),
    .S1_G_B2(\net_Lut-U178_0_S1_G_B2_to_G27_7_0 ),
    .S1_G_B3(\net_Lut-U174_0_S1_G_B3_to_G37_7_0 ),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U141_0_X_to_S1_X7_7_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U173_1_Y_to_S1_Y7_7_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_e21.CONF = "10";
  defparam GSB_CNT_7_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_h6w10.CONF = "000";
  defparam GSB_CNT_7_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_out2.CONF = "011110";
  defparam GSB_CNT_7_8_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_7_8_0_inst.sps_out4.CONF = "000111";
  defparam GSB_CNT_7_8_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_out6.CONF = "001011";
  defparam GSB_CNT_7_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s0_f_b1.CONF = "100111011";
  defparam GSB_CNT_7_8_0_inst.sps_s0_f_b2.CONF = "100111011";
  defparam GSB_CNT_7_8_0_inst.sps_s0_f_b3.CONF = "100111110";
  defparam GSB_CNT_7_8_0_inst.sps_s0_f_b4.CONF = "010111101";
  defparam GSB_CNT_7_8_0_inst.sps_s0_g_b1.CONF = "100011";
  defparam GSB_CNT_7_8_0_inst.sps_s0_g_b2.CONF = "011101";
  defparam GSB_CNT_7_8_0_inst.sps_s0_g_b3.CONF = "100101";
  defparam GSB_CNT_7_8_0_inst.sps_s0_g_b4.CONF = "110111";
  defparam GSB_CNT_7_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s16.CONF = "10";
  defparam GSB_CNT_7_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s1_f_b1.CONF = "100111101";
  defparam GSB_CNT_7_8_0_inst.sps_s1_f_b2.CONF = "011101111";
  defparam GSB_CNT_7_8_0_inst.sps_s1_f_b3.CONF = "110111111";
  defparam GSB_CNT_7_8_0_inst.sps_s1_f_b4.CONF = "100111101";
  defparam GSB_CNT_7_8_0_inst.sps_s1_g_b1.CONF = "011010";
  defparam GSB_CNT_7_8_0_inst.sps_s1_g_b2.CONF = "010000";
  defparam GSB_CNT_7_8_0_inst.sps_s1_g_b3.CONF = "010101";
  defparam GSB_CNT_7_8_0_inst.sps_s1_g_b4.CONF = "011111";
  defparam GSB_CNT_7_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_s2.CONF = "01";
  defparam GSB_CNT_7_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s4.CONF = "10";
  defparam GSB_CNT_7_8_0_inst.sps_s5.CONF = "10";
  defparam GSB_CNT_7_8_0_inst.sps_s6.CONF = "10";
  defparam GSB_CNT_7_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_v6n0.CONF = "0100";
  defparam GSB_CNT_7_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_v6n3.CONF = "0100";
  defparam GSB_CNT_7_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_v6s0.CONF = "0011";
  defparam GSB_CNT_7_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_8_0_inst.sps_v6s3.CONF = "0011";
  defparam GSB_CNT_7_8_0_inst.sps_v6s4.CONF = "011";
  defparam GSB_CNT_7_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w11.CONF = "10";
  defparam GSB_CNT_7_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w19.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e15_w15.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_e9_w9.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n18_e14.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n19_e19.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n1_w2.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s0_w2.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s10_w8.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_s11_e9.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s21_w3.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s2_e20.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s4_e2.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s9_e11.CONF = "0";
  defparam GSB_CNT_7_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_8_0_inst (
    .E0(),
    .E1(),
    .E2(\net_cnt_lcd_reg[0]_E2_to_W27_9_0 ),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(\net_Lut-U176_0_1_W7_to_E77_8_0 ),
    .E8(),
    .E9(\net_Lut-U201_0_0_W9_to_E97_8_0 ),
    .E10(),
    .E11(\net_Lut-U189_2_E11_to_W117_9_0 ),
    .E12(),
    .E13(),
    .E14(\net_cnt_lcd_reg[3]_E14_to_W147_9_0 ),
    .E15(\net_cnt_lcd_reg[7]_E15_to_W157_9_0 ),
    .E16(),
    .E17(),
    .E18(),
    .E19(\net_Lut-U201_0_0_W19_to_E197_8_0 ),
    .E20(\net_cnt_lcd_reg[1]_E20_to_W207_9_0 ),
    .E21(\net_cnt_lcd_reg[0]_E21_to_W217_9_0 ),
    .E22(),
    .E23(\net_Lut-U130_0_1_W23_to_E237_8_0 ),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(\net_cnt_lcd_reg[3]_S4_to_N47_8_0 ),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(\net_Lut-U144_0_0_S14_to_N147_8_0 ),
    .N15(),
    .N16(),
    .N17(),
    .N18(\net_cnt_lcd_reg[3]_S18_to_N187_8_0 ),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(\net_cnt_lcd_reg[5]_E2_to_W27_8_0 ),
    .W3(\net_Lut-U178_0_W3_to_E37_7_0 ),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(\net_cnt_lcd_reg[4]_E8_to_W87_8_0 ),
    .W9(\net_Lut-U201_0_0_W9_to_E97_7_0 ),
    .W10(),
    .W11(\net_Lut-U174_0_W11_to_E117_7_0 ),
    .W12(),
    .W13(),
    .W14(\net_cnt_lcd_reg[6]_E14_to_W147_8_0 ),
    .W15(\net_cnt_lcd_reg[7]_E15_to_W157_8_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(\net_Lut-U138_0_W19_to_E197_7_0 ),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(\net_cnt_lcd_reg[1]_S2_to_N28_8_0 ),
    .S3(),
    .S4(\net_cnt_lcd_reg[0]_S4_to_N48_8_0 ),
    .S5(),
    .S6(\net_cnt_lcd_reg[1]_S6_to_N68_8_0 ),
    .S7(),
    .S8(),
    .S9(\net_Lut-U189_2_N9_to_S97_8_0 ),
    .S10(),
    .S11(\net_Lut-U201_0_0_S11_to_N118_8_0 ),
    .S12(),
    .S13(),
    .S14(\net_Lut-U209_0_0_N14_to_S147_8_0 ),
    .S15(),
    .S16(\net_Lut-U232_0_0_S16_to_N168_8_0 ),
    .S17(\net_Lut-U204_0_1_N17_to_S177_8_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(\net_Lut-U178_0_N21_to_S217_8_0 ),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(\net_cnt_lcd_reg[1]_H6E0_to_H6M07_8_0 ),
    .H6M1(),
    .H6M2(),
    .H6M3(\net_cnt_lcd_reg[0]_H6E3_to_H6M37_8_0 ),
    .H6M4(),
    .H6M5(\net_cnt_lcd_reg[0]_H6E5_to_H6M57_8_0 ),
    .H6M6(),
    .H6M7(\net_Lut-U232_0_0_H6E7_to_H6M77_8_0 ),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(\net_Lut-U126_1_H6W10_to_LEFT_H6E107_2_0 ),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(\net_Lut-U175_0_0_OUT0_to_OUT_W07_8_0 ),
    .OUT_W1(),
    .OUT_E6(\net_Lut-U127_0_OUT6_to_OUT_E67_8_0 ),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(\net_cnt_lcd_reg[1]_V6S0_to_V6M010_8_0 ),
    .V6S1(),
    .V6S2(),
    .V6S3(\net_cnt_lcd_reg[0]_V6S3_to_V6M310_8_0 ),
    .V6S4(\net_cnt_lcd_reg[0]_V6S4_to_V6M410_8_0 ),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U144_0_0_S0_F_B1_to_F17_8_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[4]_S0_F_B2_to_F27_8_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[5]_S0_F_B3_to_F37_8_0 ),
    .S0_F_B4(\net_cnt_lcd_reg[6]_S0_F_B4_to_F47_8_0 ),
    .S0_G_B1(\net_Lut-U126_0_0_S0_G_B1_to_G17_8_0 ),
    .S0_G_B2(\net_Lut-U130_0_1_S0_G_B2_to_G27_8_0 ),
    .S0_G_B3(\net_Lut-U209_0_0_S0_G_B3_to_G37_8_0 ),
    .S0_G_B4(\net_Lut-U127_0_S0_G_B4_to_G47_8_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U138_0_X_to_S0_X7_8_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U126_1_Y_to_S0_Y7_8_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U232_0_0_S1_F_B1_to_F17_8_0 ),
    .S1_F_B2(\net_Lut-U176_0_1_S1_F_B2_to_F27_8_0 ),
    .S1_F_B3(\net_Lut-U175_0_0_S1_F_B3_to_F37_8_0 ),
    .S1_F_B4(\net_Lut-U204_0_1_S1_F_B4_to_F47_8_0 ),
    .S1_G_B1(\net_cnt_lcd_reg[5]_S1_G_B1_to_G17_8_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[3]_S1_G_B2_to_G27_8_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[4]_S1_G_B3_to_G37_8_0 ),
    .S1_G_B4(\net_Lut-U201_0_0_S1_G_B4_to_G47_8_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U174_0_X_to_S1_X7_8_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U126_0_0_Y_to_S1_Y7_8_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e3.CONF = "10";
  defparam GSB_CNT_8_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e5.CONF = "10";
  defparam GSB_CNT_8_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_6_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_n6.CONF = "10";
  defparam GSB_CNT_8_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_n9.CONF = "10";
  defparam GSB_CNT_8_6_0_inst.sps_out0.CONF = "011110";
  defparam GSB_CNT_8_6_0_inst.sps_out1.CONF = "011101";
  defparam GSB_CNT_8_6_0_inst.sps_out2.CONF = "000111";
  defparam GSB_CNT_8_6_0_inst.sps_out3.CONF = "001011";
  defparam GSB_CNT_8_6_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_f_b1.CONF = "100111101";
  defparam GSB_CNT_8_6_0_inst.sps_s0_f_b2.CONF = "001111101";
  defparam GSB_CNT_8_6_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_g_b1.CONF = "100101";
  defparam GSB_CNT_8_6_0_inst.sps_s0_g_b2.CONF = "010101";
  defparam GSB_CNT_8_6_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_f_b1.CONF = "100011111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_f_b2.CONF = "011111110";
  defparam GSB_CNT_8_6_0_inst.sps_s1_f_b3.CONF = "010011111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_g_b1.CONF = "100100";
  defparam GSB_CNT_8_6_0_inst.sps_s1_g_b2.CONF = "100111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_g_b3.CONF = "001111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s0.CONF = "0000";
  defparam GSB_CNT_8_6_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e18_w18.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_e19_w19.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n12_e8.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n13_e13.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n15_e15.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n17_e17.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n1_e1.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n4_e0.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n7_e7.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s0_n0.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s11_e9.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s12_n12.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s16_w18.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s1_n1.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s22_w20.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s23_e21.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s2_n2.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s3_n3.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s5_n5.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s7_n7.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s9_e11.CONF = "0";
  defparam GSB_CNT_8_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_6_0_inst (
    .E0(net_U113_W0_to_E08_6_0),
    .E1(\net_cnt_lcd_reg[5]_E1_to_W18_7_0 ),
    .E2(),
    .E3(\net_Lut-U190_0_1_E3_to_W38_7_0 ),
    .E4(),
    .E5(\net_Lut-U190_0_1_E5_to_W58_7_0 ),
    .E6(),
    .E7(\net_cnt_lcd_reg[4]_E7_to_W78_7_0 ),
    .E8(\net_cnt_lcd_reg[7]_E8_to_W88_7_0 ),
    .E9(\net_Lut-U191_1_W9_to_E98_6_0 ),
    .E10(),
    .E11(),
    .E12(),
    .E13(\net_cnt_lcd_reg[6]_E13_to_W138_7_0 ),
    .E14(),
    .E15(net_U113_W15_to_E158_6_0),
    .E16(),
    .E17(\net_cnt_lcd_reg[5]_E17_to_W178_7_0 ),
    .E18(\net_cnt_lcd_reg[0]_E18_to_W188_7_0 ),
    .E19(\net_Lut-U232_0_0_E19_to_W198_7_0 ),
    .E20(),
    .E21(\net_Lut-U137_0_0_W21_to_E218_6_0 ),
    .E22(),
    .E23(),
    .N0(\net_cnt_lcd_reg[5]_S0_to_N08_6_0 ),
    .N1(\net_cnt_lcd_reg[5]_S1_to_N18_6_0 ),
    .N2(\net_cnt_lcd_reg[5]_S2_to_N28_6_0 ),
    .N3(\net_cnt_lcd_reg[1]_S3_to_N38_6_0 ),
    .N4(net_U113_N4_to_S47_6_0),
    .N5(\net_cnt_lcd_reg[4]_S5_to_N58_6_0 ),
    .N6(\net_Lut-U143_0_N6_to_S67_6_0 ),
    .N7(\net_cnt_lcd_reg[4]_S7_to_N78_6_0 ),
    .N8(),
    .N9(\net_Lut-U136_0_N9_to_S97_6_0 ),
    .N10(),
    .N11(),
    .N12(\net_cnt_lcd_reg[7]_S12_to_N128_6_0 ),
    .N13(\net_cnt_lcd_reg[6]_S13_to_N138_6_0 ),
    .N14(\net_cnt_lcd_reg[7]_S14_to_N148_6_0 ),
    .N15(net_U113_N15_to_S157_6_0),
    .N16(),
    .N17(\net_cnt_lcd_reg[5]_S17_to_N178_6_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_cnt_lcd_reg[3]_E12_to_W128_6_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(\net_cnt_lcd_reg[0]_E18_to_W188_6_0 ),
    .W19(\net_Lut-U232_0_0_E19_to_W198_6_0 ),
    .W20(\net_cnt_lcd_reg[1]_E20_to_W208_6_0 ),
    .W21(),
    .W22(),
    .W23(),
    .S0(\net_cnt_lcd_reg[5]_S0_to_N09_6_0 ),
    .S1(\net_cnt_lcd_reg[5]_S1_to_N19_6_0 ),
    .S2(\net_cnt_lcd_reg[5]_S2_to_N29_6_0 ),
    .S3(\net_cnt_lcd_reg[1]_S3_to_N39_6_0 ),
    .S4(),
    .S5(\net_cnt_lcd_reg[4]_S5_to_N59_6_0 ),
    .S6(),
    .S7(\net_cnt_lcd_reg[4]_S7_to_N79_6_0 ),
    .S8(),
    .S9(\net_Lut-U144_0_0_N9_to_S98_6_0 ),
    .S10(),
    .S11(\net_Lut-U191_1_S11_to_N119_6_0 ),
    .S12(\net_cnt_lcd_reg[7]_S12_to_N129_6_0 ),
    .S13(),
    .S14(),
    .S15(),
    .S16(\net_cnt_lcd_reg[0]_S16_to_N169_6_0 ),
    .S17(),
    .S18(),
    .S19(),
    .S20(\net_cnt_lcd_reg[3]_N20_to_S208_6_0 ),
    .S21(),
    .S22(\net_cnt_lcd_reg[1]_S22_to_N229_6_0 ),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(\net_Lut-U186_0_V6S0_to_V6M011_6_0 ),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[4]_S0_F_B1_to_F18_6_0 ),
    .S0_F_B2(\net_Lut-U144_0_0_S0_F_B2_to_F28_6_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_cnt_lcd_reg[7]_S0_G_B1_to_G18_6_0 ),
    .S0_G_B2(\net_Lut-U137_0_0_S0_G_B2_to_G28_6_0 ),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U143_0_X_to_S0_X8_6_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U136_0_Y_to_S0_Y8_6_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[1]_S1_F_B1_to_F18_6_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[3]_S1_F_B2_to_F28_6_0 ),
    .S1_F_B3(\net_cnt_lcd_reg[5]_S1_F_B3_to_F38_6_0 ),
    .S1_F_B4(),
    .S1_G_B1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G18_6_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[5]_S1_G_B2_to_G28_6_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[3]_S1_G_B3_to_G38_6_0 ),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U190_0_1_X_to_S1_X8_6_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U186_0_Y_to_S1_Y8_6_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_7_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_e17.CONF = "10";
  defparam GSB_CNT_8_7_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_e21.CONF = "10";
  defparam GSB_CNT_8_7_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_7_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_7_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n13.CONF = "10";
  defparam GSB_CNT_8_7_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_n9.CONF = "10";
  defparam GSB_CNT_8_7_0_inst.sps_out0.CONF = "011110";
  defparam GSB_CNT_8_7_0_inst.sps_out1.CONF = "011110";
  defparam GSB_CNT_8_7_0_inst.sps_out2.CONF = "001011";
  defparam GSB_CNT_8_7_0_inst.sps_out3.CONF = "001011";
  defparam GSB_CNT_8_7_0_inst.sps_out4.CONF = "011101";
  defparam GSB_CNT_8_7_0_inst.sps_out5.CONF = "011110";
  defparam GSB_CNT_8_7_0_inst.sps_out6.CONF = "000111";
  defparam GSB_CNT_8_7_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s0_f_b1.CONF = "010111110";
  defparam GSB_CNT_8_7_0_inst.sps_s0_f_b2.CONF = "100111011";
  defparam GSB_CNT_8_7_0_inst.sps_s0_f_b3.CONF = "001111011";
  defparam GSB_CNT_8_7_0_inst.sps_s0_f_b4.CONF = "010111011";
  defparam GSB_CNT_8_7_0_inst.sps_s0_g_b1.CONF = "010100";
  defparam GSB_CNT_8_7_0_inst.sps_s0_g_b2.CONF = "100000";
  defparam GSB_CNT_8_7_0_inst.sps_s0_g_b3.CONF = "011011";
  defparam GSB_CNT_8_7_0_inst.sps_s0_g_b4.CONF = "010000";
  defparam GSB_CNT_8_7_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s1_f_b1.CONF = "010111011";
  defparam GSB_CNT_8_7_0_inst.sps_s1_f_b2.CONF = "100011111";
  defparam GSB_CNT_8_7_0_inst.sps_s1_f_b3.CONF = "010101111";
  defparam GSB_CNT_8_7_0_inst.sps_s1_f_b4.CONF = "100101111";
  defparam GSB_CNT_8_7_0_inst.sps_s1_g_b1.CONF = "010101";
  defparam GSB_CNT_8_7_0_inst.sps_s1_g_b2.CONF = "100100";
  defparam GSB_CNT_8_7_0_inst.sps_s1_g_b3.CONF = "100100";
  defparam GSB_CNT_8_7_0_inst.sps_s1_g_b4.CONF = "011101";
  defparam GSB_CNT_8_7_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_s2.CONF = "01";
  defparam GSB_CNT_8_7_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_7_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_v6n0.CONF = "0001";
  defparam GSB_CNT_8_7_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_v6n3.CONF = "0100";
  defparam GSB_CNT_8_7_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_7_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_7_0_inst.sps_w0.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_w15.CONF = "10";
  defparam GSB_CNT_8_7_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w21.CONF = "10";
  defparam GSB_CNT_8_7_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_7_0_inst.sps_w9.CONF = "10";
  defparam GSB_CNT_8_7_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e13_w13.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e1_w1.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e5_w5.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e7_w7.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n15_e15.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n18_e14.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n23_e23.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s10_n10.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s11_w13.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s21_w3.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s5_n5.CONF = "0";
  defparam GSB_CNT_8_7_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_7_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_7_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(\net_Lut-U190_0_1_E5_to_W58_8_0 ),
    .E6(),
    .E7(\net_cnt_lcd_reg[4]_E7_to_W78_8_0 ),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(\net_Lut-U225_0_E14_to_W148_8_0 ),
    .E15(\net_cnt_lcd_reg[7]_E15_to_W158_8_0 ),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(\net_Lut-U188_0_0_E21_to_W218_8_0 ),
    .E22(),
    .E23(\net_cnt_lcd_reg[3]_W23_to_E238_7_0 ),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(\net_Lut-U205_0_0_S5_to_N58_7_0 ),
    .N6(),
    .N7(),
    .N8(),
    .N9(\net_Lut-U191_1_N9_to_S97_7_0 ),
    .N10(\net_cnt_lcd_reg[4]_S10_to_N108_7_0 ),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(\net_cnt_lcd_reg[7]_S15_to_N158_7_0 ),
    .N16(),
    .N17(),
    .N18(\net_Lut-U225_0_S18_to_N188_7_0 ),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(net_U113_W0_to_E08_6_0),
    .W1(\net_cnt_lcd_reg[5]_E1_to_W18_7_0 ),
    .W2(),
    .W3(\net_Lut-U190_0_1_E3_to_W38_7_0 ),
    .W4(),
    .W5(\net_Lut-U190_0_1_E5_to_W58_7_0 ),
    .W6(),
    .W7(\net_cnt_lcd_reg[4]_E7_to_W78_7_0 ),
    .W8(\net_cnt_lcd_reg[7]_E8_to_W88_7_0 ),
    .W9(\net_Lut-U191_1_W9_to_E98_6_0 ),
    .W10(),
    .W11(),
    .W12(),
    .W13(\net_cnt_lcd_reg[6]_E13_to_W138_7_0 ),
    .W14(),
    .W15(net_U113_W15_to_E158_6_0),
    .W16(),
    .W17(\net_cnt_lcd_reg[5]_E17_to_W178_7_0 ),
    .W18(\net_cnt_lcd_reg[0]_E18_to_W188_7_0 ),
    .W19(\net_Lut-U232_0_0_E19_to_W198_7_0 ),
    .W20(),
    .W21(\net_Lut-U137_0_0_W21_to_E218_6_0 ),
    .W22(),
    .W23(),
    .S0(),
    .S1(\net_cnt_lcd_reg[2]_N1_to_S18_7_0 ),
    .S2(\net_Lut-U213_0_0_S2_to_N29_7_0 ),
    .S3(),
    .S4(),
    .S5(\net_Lut-U205_0_0_S5_to_N59_7_0 ),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(\net_Lut-U144_0_0_N12_to_S128_7_0 ),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(\net_Lut-U190_0_1_S21_to_N219_7_0 ),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(\net_Lut-U188_0_0_H6W3_to_H6M38_7_0 ),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(\net_Lut-U213_0_0_OUT1_to_OUT_W18_8_0 ),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(net_U113_V6N2_to_V6M28_7_0),
    .V6M3(),
    .V6M4(),
    .V6M5(net_U113_V6N5_to_V6M58_7_0),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U144_0_0_S0_F_B1_to_F18_7_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[4]_S0_F_B2_to_F28_7_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[5]_S0_F_B3_to_F38_7_0 ),
    .S0_F_B4(\net_cnt_lcd_reg[6]_S0_F_B4_to_F48_7_0 ),
    .S0_G_B1(\net_cnt_lcd_reg[3]_S0_G_B1_to_G18_7_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[2]_S0_G_B2_to_G28_7_0 ),
    .S0_G_B3(\net_Lut-U193_0_0_S0_G_B3_to_G38_7_0 ),
    .S0_G_B4(\net_Lut-U213_0_0_S0_G_B4_to_G48_7_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U137_0_0_X_to_S0_X8_7_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U191_1_Y_to_S0_Y8_7_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[4]_S1_F_B1_to_F18_7_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[7]_S1_F_B2_to_F28_7_0 ),
    .S1_F_B3(\net_Lut-U232_0_0_S1_F_B3_to_F38_7_0 ),
    .S1_F_B4(\net_cnt_lcd_reg[5]_S1_F_B4_to_F48_7_0 ),
    .S1_G_B1(\net_cnt_lcd_reg[4]_S1_G_B1_to_G18_7_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[7]_S1_G_B2_to_G28_7_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[6]_S1_G_B3_to_G38_7_0 ),
    .S1_G_B4(\net_cnt_lcd_reg[0]_S1_G_B4_to_G48_7_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U193_0_0_X_to_S1_X8_7_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U213_0_0_Y_to_S1_Y8_7_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_9_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_h6w1.CONF = "0010";
  defparam GSB_CNT_8_9_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_9_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_9_0_inst.sps_n0.CONF = "01";
  defparam GSB_CNT_8_9_0_inst.sps_n1.CONF = "10";
  defparam GSB_CNT_8_9_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_out0.CONF = "000111";
  defparam GSB_CNT_8_9_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_out2.CONF = "011110";
  defparam GSB_CNT_8_9_0_inst.sps_out3.CONF = "001011";
  defparam GSB_CNT_8_9_0_inst.sps_out4.CONF = "000111";
  defparam GSB_CNT_8_9_0_inst.sps_out5.CONF = "001011";
  defparam GSB_CNT_8_9_0_inst.sps_out6.CONF = "011101";
  defparam GSB_CNT_8_9_0_inst.sps_out7.CONF = "001011";
  defparam GSB_CNT_8_9_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_s0_f_b1.CONF = "100111101";
  defparam GSB_CNT_8_9_0_inst.sps_s0_f_b2.CONF = "100110111";
  defparam GSB_CNT_8_9_0_inst.sps_s0_f_b3.CONF = "001111110";
  defparam GSB_CNT_8_9_0_inst.sps_s0_f_b4.CONF = "010011111";
  defparam GSB_CNT_8_9_0_inst.sps_s0_g_b1.CONF = "011100";
  defparam GSB_CNT_8_9_0_inst.sps_s0_g_b2.CONF = "011011";
  defparam GSB_CNT_8_9_0_inst.sps_s0_g_b3.CONF = "010000";
  defparam GSB_CNT_8_9_0_inst.sps_s0_g_b4.CONF = "100011";
  defparam GSB_CNT_8_9_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_s13.CONF = "10";
  defparam GSB_CNT_8_9_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_s1_f_b1.CONF = "001110111";
  defparam GSB_CNT_8_9_0_inst.sps_s1_f_b2.CONF = "010111110";
  defparam GSB_CNT_8_9_0_inst.sps_s1_f_b3.CONF = "010101111";
  defparam GSB_CNT_8_9_0_inst.sps_s1_f_b4.CONF = "100111011";
  defparam GSB_CNT_8_9_0_inst.sps_s1_g_b1.CONF = "001111";
  defparam GSB_CNT_8_9_0_inst.sps_s1_g_b2.CONF = "010000";
  defparam GSB_CNT_8_9_0_inst.sps_s1_g_b3.CONF = "011011";
  defparam GSB_CNT_8_9_0_inst.sps_s1_g_b4.CONF = "100101";
  defparam GSB_CNT_8_9_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s5.CONF = "10";
  defparam GSB_CNT_8_9_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_s8.CONF = "01";
  defparam GSB_CNT_8_9_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_9_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_v6s10.CONF = "001";
  defparam GSB_CNT_8_9_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_9_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_9_0_inst.sps_v6s8.CONF = "001";
  defparam GSB_CNT_8_9_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w17.CONF = "10";
  defparam GSB_CNT_8_9_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w6.CONF = "01";
  defparam GSB_CNT_8_9_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_9_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e19_w19.CONF = "0";
  defparam GSB_CNT_8_9_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n4_e0.CONF = "0";
  defparam GSB_CNT_8_9_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n6_e2.CONF = "0";
  defparam GSB_CNT_8_9_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_n9_w10.CONF = "0";
  defparam GSB_CNT_8_9_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s17_n17.CONF = "0";
  defparam GSB_CNT_8_9_0_inst.switch_s17_w23.CONF = "0";
  defparam GSB_CNT_8_9_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s22_e16.CONF = "0";
  defparam GSB_CNT_8_9_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s2_w0.CONF = "0";
  defparam GSB_CNT_8_9_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_9_0_inst.switch_s9_n9.CONF = "0";
  defparam GSB_CNT_8_9_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_9_0_inst (
    .E0(\net_cnt_lcd_reg[5]_E0_to_W08_10_0 ),
    .E1(),
    .E2(\net_cnt_lcd_reg[5]_E2_to_W28_10_0 ),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(\net_Lut-U229_0_W16_to_E168_9_0 ),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(\net_Lut-U176_0_1_N0_to_S07_9_0 ),
    .N1(\net_Lut-U176_0_1_N1_to_S17_9_0 ),
    .N2(),
    .N3(),
    .N4(\net_cnt_lcd_reg[5]_S4_to_N48_9_0 ),
    .N5(),
    .N6(\net_cnt_lcd_reg[5]_S6_to_N68_9_0 ),
    .N7(),
    .N8(),
    .N9(\net_cnt_lcd_reg[4]_S9_to_N98_9_0 ),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(\net_cnt_lcd_reg[6]_S17_to_N178_9_0 ),
    .N18(\net_cnt_lcd_reg[7]_S18_to_N188_9_0 ),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(\net_cnt_lcd_reg[0]_E0_to_W08_9_0 ),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(\net_Lut-U202_0_0_W6_to_E68_8_0 ),
    .W7(\net_cnt_lcd_reg[2]_E7_to_W78_9_0 ),
    .W8(),
    .W9(),
    .W10(\net_cnt_lcd_reg[4]_W10_to_E108_8_0 ),
    .W11(\net_cnt_lcd_reg[1]_E11_to_W118_9_0 ),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(\net_Lut-U204_0_1_W17_to_E178_8_0 ),
    .W18(),
    .W19(\net_cnt_lcd_reg[3]_E19_to_W198_9_0 ),
    .W20(),
    .W21(),
    .W22(\net_cnt_lcd_reg[1]_E22_to_W228_9_0 ),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(\net_Lut-U204_0_1_S8_to_N89_9_0 ),
    .S9(\net_cnt_lcd_reg[4]_S9_to_N99_9_0 ),
    .S10(),
    .S11(),
    .S12(),
    .S13(\net_Lut-U176_0_1_S13_to_N139_9_0 ),
    .S14(),
    .S15(),
    .S16(),
    .S17(\net_cnt_lcd_reg[6]_S17_to_N179_9_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(\net_Lut-U229_0_S22_to_N229_9_0 ),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(\net_Lut-U180_0_0_OUT6_to_OUT_E68_8_0 ),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(\net_Lut-U202_0_0_V6N9_to_V6M98_9_0 ),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(\net_Lut-U204_0_1_V6S8_to_V6M811_9_0 ),
    .V6S9(),
    .V6S10(\net_Lut-U204_0_1_V6S10_to_V6M1011_9_0 ),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U176_0_0_S0_F_B1_to_F18_9_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[7]_S0_F_B2_to_F28_9_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[6]_S0_F_B3_to_F38_9_0 ),
    .S0_F_B4(\net_cnt_lcd_reg[0]_S0_F_B4_to_F48_9_0 ),
    .S0_G_B1(\net_cnt_lcd_reg[1]_S0_G_B1_to_G18_9_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[4]_S0_G_B2_to_G28_9_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[5]_S0_G_B3_to_G38_9_0 ),
    .S0_G_B4(\net_cnt_lcd_reg[3]_S0_G_B4_to_G48_9_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U176_0_1_X_to_S0_X8_9_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U204_0_1_Y_to_S0_Y8_9_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[1]_S1_F_B1_to_F18_9_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[5]_S1_F_B2_to_F28_9_0 ),
    .S1_F_B3(\net_cnt_lcd_reg[3]_S1_F_B3_to_F38_9_0 ),
    .S1_F_B4(\net_cnt_lcd_reg[2]_S1_F_B4_to_F48_9_0 ),
    .S1_G_B1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G18_9_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[5]_S1_G_B2_to_G28_9_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[4]_S1_G_B3_to_G38_9_0 ),
    .S1_G_B4(\net_cnt_lcd_reg[2]_S1_G_B4_to_G48_9_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U180_0_0_X_to_S1_X8_9_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U176_0_0_Y_to_S1_Y8_9_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_10_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_h6w2.CONF = "0011";
  defparam GSB_CNT_7_10_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_10_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_10_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n21.CONF = "10";
  defparam GSB_CNT_7_10_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_out2.CONF = "011101";
  defparam GSB_CNT_7_10_0_inst.sps_out3.CONF = "001011";
  defparam GSB_CNT_7_10_0_inst.sps_out4.CONF = "011101";
  defparam GSB_CNT_7_10_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_out6.CONF = "011110";
  defparam GSB_CNT_7_10_0_inst.sps_out7.CONF = "000111";
  defparam GSB_CNT_7_10_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_s0_f_b1.CONF = "100111110";
  defparam GSB_CNT_7_10_0_inst.sps_s0_f_b2.CONF = "100110111";
  defparam GSB_CNT_7_10_0_inst.sps_s0_f_b3.CONF = "001111110";
  defparam GSB_CNT_7_10_0_inst.sps_s0_f_b4.CONF = "100111011";
  defparam GSB_CNT_7_10_0_inst.sps_s0_g_b1.CONF = "001010";
  defparam GSB_CNT_7_10_0_inst.sps_s0_g_b2.CONF = "100011";
  defparam GSB_CNT_7_10_0_inst.sps_s0_g_b3.CONF = "011010";
  defparam GSB_CNT_7_10_0_inst.sps_s0_g_b4.CONF = "011010";
  defparam GSB_CNT_7_10_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s15.CONF = "10";
  defparam GSB_CNT_7_10_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_s1_f_b1.CONF = "100111110";
  defparam GSB_CNT_7_10_0_inst.sps_s1_f_b2.CONF = "011110111";
  defparam GSB_CNT_7_10_0_inst.sps_s1_f_b3.CONF = "100110111";
  defparam GSB_CNT_7_10_0_inst.sps_s1_f_b4.CONF = "100011111";
  defparam GSB_CNT_7_10_0_inst.sps_s1_g_b1.CONF = "011000";
  defparam GSB_CNT_7_10_0_inst.sps_s1_g_b2.CONF = "001010";
  defparam GSB_CNT_7_10_0_inst.sps_s1_g_b3.CONF = "010111";
  defparam GSB_CNT_7_10_0_inst.sps_s1_g_b4.CONF = "010000";
  defparam GSB_CNT_7_10_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s5.CONF = "10";
  defparam GSB_CNT_7_10_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_10_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_10_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_7_10_0_inst.sps_v6s8.CONF = "001";
  defparam GSB_CNT_7_10_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w19.CONF = "0";
  defparam GSB_CNT_7_10_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_10_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e5_w5.CONF = "0";
  defparam GSB_CNT_7_10_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n11_w12.CONF = "0";
  defparam GSB_CNT_7_10_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n12_w17.CONF = "0";
  defparam GSB_CNT_7_10_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n1_w2.CONF = "0";
  defparam GSB_CNT_7_10_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s7_e5.CONF = "0";
  defparam GSB_CNT_7_10_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_10_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_10_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(\net_cnt_lcd_reg[1]_W5_to_E57_10_0 ),
    .E6(\net_cnt_lcd_reg[1]_W6_to_E67_10_0 ),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(\net_cnt_lcd_reg[0]_W20_to_E207_10_0 ),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(\net_cnt_lcd_reg[3]_S8_to_N87_10_0 ),
    .N9(),
    .N10(\net_cnt_lcd_reg[2]_S10_to_N107_10_0 ),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(\net_cnt_lcd_reg[3]_S18_to_N187_10_0 ),
    .N19(),
    .N20(),
    .N21(),
    .N22(\net_cnt_lcd_reg[2]_S22_to_N227_10_0 ),
    .N23(),
    .W0(),
    .W1(),
    .W2(\net_cnt_lcd_reg[5]_E2_to_W27_10_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(\net_cnt_lcd_reg[4]_E6_to_W67_10_0 ),
    .W7(),
    .W8(),
    .W9(\net_cnt_lcd_reg[4]_E9_to_W97_10_0 ),
    .W10(),
    .W11(),
    .W12(\net_cnt_lcd_reg[7]_E12_to_W127_10_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(\net_cnt_lcd_reg[6]_E17_to_W177_10_0 ),
    .W18(),
    .W19(\net_Lut-U229_0_W19_to_E197_9_0 ),
    .W20(),
    .W21(),
    .W22(),
    .W23(\net_cnt_lcd_reg[5]_E23_to_W237_10_0 ),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(\net_Lut-U229_0_S5_to_N58_10_0 ),
    .S6(),
    .S7(\net_cnt_lcd_reg[1]_S7_to_N78_10_0 ),
    .S8(),
    .S9(\net_Lut-U177_0_0_N9_to_S97_10_0 ),
    .S10(),
    .S11(),
    .S12(\net_Lut-U183_0_0_N12_to_S127_10_0 ),
    .S13(),
    .S14(),
    .S15(\net_Lut-U229_0_S15_to_N158_10_0 ),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(\net_Lut-U225_0_H6W2_to_H6M27_7_0 ),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(\net_Lut-U127_0_0_OUT6_to_OUT_E67_9_0 ),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(\net_Lut-U225_0_V6N2_to_V6M27_10_0 ),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(\net_Lut-U154_0_V6S8_to_V6M810_10_0 ),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[1]_S0_F_B1_to_F17_10_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[3]_S0_F_B2_to_F27_10_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[5]_S0_F_B3_to_F37_10_0 ),
    .S0_F_B4(\net_cnt_lcd_reg[2]_S0_F_B4_to_F47_10_0 ),
    .S0_G_B1(\net_cnt_lcd_reg[2]_S0_G_B1_to_G17_10_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G27_10_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[3]_S0_G_B3_to_G37_10_0 ),
    .S0_G_B4(\net_cnt_lcd_reg[5]_S0_G_B4_to_G47_10_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U129_0_X_to_S0_X7_10_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U154_0_Y_to_S0_Y7_10_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[4]_S1_F_B1_to_F17_10_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[7]_S1_F_B2_to_F27_10_0 ),
    .S1_F_B3(\net_cnt_lcd_reg[6]_S1_F_B3_to_F37_10_0 ),
    .S1_F_B4(\net_cnt_lcd_reg[0]_S1_F_B4_to_F47_10_0 ),
    .S1_G_B1(\net_Lut-U177_0_0_S1_G_B1_to_G17_10_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[4]_S1_G_B2_to_G27_10_0 ),
    .S1_G_B3(\net_Lut-U129_0_S1_G_B3_to_G37_10_0 ),
    .S1_G_B4(\net_Lut-U183_0_0_S1_G_B4_to_G47_10_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U229_0_X_to_S1_X7_10_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U127_0_0_Y_to_S1_Y7_10_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_9_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_e0.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e12.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_e21.CONF = "01";
  defparam GSB_CNT_10_9_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_e7.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.sps_e8.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_9_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_9_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n1.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_n16.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.sps_n17.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n23.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n5.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_n9.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.sps_out0.CONF = "000111";
  defparam GSB_CNT_10_9_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_out2.CONF = "011110";
  defparam GSB_CNT_10_9_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_10_9_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_out5.CONF = "001011";
  defparam GSB_CNT_10_9_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s0_f_b1.CONF = "010011111";
  defparam GSB_CNT_10_9_0_inst.sps_s0_f_b2.CONF = "010101111";
  defparam GSB_CNT_10_9_0_inst.sps_s0_f_b3.CONF = "010111101";
  defparam GSB_CNT_10_9_0_inst.sps_s0_f_b4.CONF = "110111111";
  defparam GSB_CNT_10_9_0_inst.sps_s0_g_b1.CONF = "010100";
  defparam GSB_CNT_10_9_0_inst.sps_s0_g_b2.CONF = "010010";
  defparam GSB_CNT_10_9_0_inst.sps_s0_g_b3.CONF = "010011";
  defparam GSB_CNT_10_9_0_inst.sps_s0_g_b4.CONF = "001101";
  defparam GSB_CNT_10_9_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_s12.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_s16.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s1_f_b1.CONF = "100111011";
  defparam GSB_CNT_10_9_0_inst.sps_s1_f_b2.CONF = "011110111";
  defparam GSB_CNT_10_9_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_9_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_9_0_inst.sps_s1_g_b1.CONF = "100010";
  defparam GSB_CNT_10_9_0_inst.sps_s1_g_b2.CONF = "011111";
  defparam GSB_CNT_10_9_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_s2.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.sps_s20.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.sps_s21.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_s4.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_s6.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_s8.CONF = "01";
  defparam GSB_CNT_10_9_0_inst.sps_s9.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_9_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_9_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_9_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_w13.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w3.CONF = "01";
  defparam GSB_CNT_10_9_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_9_0_inst.sps_w9.CONF = "10";
  defparam GSB_CNT_10_9_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e22_w22.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e7_w7.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n11_w12.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n13_e13.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n14_w19.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n15_w16.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s15_n15.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s16_e14.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s8_w10.CONF = "0";
  defparam GSB_CNT_10_9_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_9_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_9_0_inst (
    .E0(\net_cnt_lcd_reg[5]_E0_to_W010_10_0 ),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(\net_Lut-U227_0_E8_to_W810_10_0 ),
    .E9(),
    .E10(),
    .E11(),
    .E12(\net_cnt_lcd_reg[6]_E12_to_W1210_10_0 ),
    .E13(\net_Lut-U154_0_W13_to_E1310_9_0 ),
    .E14(\net_cnt_lcd_reg[7]_E14_to_W1410_10_0 ),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(\net_cnt_lcd_reg[5]_E21_to_W2110_10_0 ),
    .E22(\net_Lut-U195_0_W22_to_E2210_9_0 ),
    .E23(),
    .N0(),
    .N1(\net_Lut-U152_0_0_N1_to_S19_9_0 ),
    .N2(),
    .N3(),
    .N4(),
    .N5(\net_cnt_lcd_reg[5]_N5_to_S59_9_0 ),
    .N6(),
    .N7(),
    .N8(),
    .N9(\net_Lut-U227_0_N9_to_S99_9_0 ),
    .N10(),
    .N11(),
    .N12(),
    .N13(\net_Lut-U154_0_N13_to_S139_9_0 ),
    .N14(\net_cnt_lcd_reg[0]_N14_to_S149_9_0 ),
    .N15(\net_Lut-U230_0_0_S15_to_N1510_9_0 ),
    .N16(),
    .N17(\net_cnt_lcd_reg[7]_N17_to_S179_9_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(\net_cnt_lcd_reg[0]_E0_to_W010_9_0 ),
    .W1(\net_cnt_lcd_reg[1]_E1_to_W110_9_0 ),
    .W2(),
    .W3(\net_Lut-U201_0_0_W3_to_E310_8_0 ),
    .W4(),
    .W5(),
    .W6(),
    .W7(\net_Lut-U201_0_0_W7_to_E710_8_0 ),
    .W8(),
    .W9(\net_Lut-U161_0_0_W9_to_E910_8_0 ),
    .W10(\net_cnt_lcd_reg[4]_W10_to_E1010_8_0 ),
    .W11(),
    .W12(\net_cnt_lcd_reg[3]_E12_to_W1210_9_0 ),
    .W13(\net_Lut-U201_0_0_W13_to_E1310_8_0 ),
    .W14(),
    .W15(),
    .W16(\net_Lut-U230_0_0_W16_to_E1610_8_0 ),
    .W17(),
    .W18(),
    .W19(\net_cnt_lcd_reg[0]_E19_to_W1910_9_0 ),
    .W20(),
    .W21(),
    .W22(\net_Lut-U195_0_W22_to_E2210_8_0 ),
    .W23(),
    .S0(),
    .S1(),
    .S2(\net_cnt_lcd_reg[4]_S2_to_N211_9_0 ),
    .S3(),
    .S4(\net_cnt_lcd_reg[5]_S4_to_N411_9_0 ),
    .S5(),
    .S6(\net_cnt_lcd_reg[5]_S6_to_N611_9_0 ),
    .S7(),
    .S8(),
    .S9(\net_cnt_lcd_reg[4]_S9_to_N911_9_0 ),
    .S10(),
    .S11(),
    .S12(\net_Lut-U170_0_S12_to_N1211_9_0 ),
    .S13(),
    .S14(),
    .S15(\net_Lut-U230_0_0_S15_to_N1511_9_0 ),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(\net_cnt_lcd_reg[7]_S20_to_N2011_9_0 ),
    .S21(\net_cnt_lcd_reg[5]_S21_to_N2111_9_0 ),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(\net_cnt_lcd_reg[5]_H6E0_to_H6M010_9_0 ),
    .H6M1(\net_cnt_lcd_reg[4]_H6W1_to_H6M110_9_0 ),
    .H6M2(\net_cnt_lcd_reg[6]_H6E2_to_H6M210_9_0 ),
    .H6M3(\net_cnt_lcd_reg[5]_H6E3_to_H6M310_9_0 ),
    .H6M4(\net_cnt_lcd_reg[4]_H6W4_to_H6M410_9_0 ),
    .H6M5(\net_cnt_lcd_reg[5]_H6E5_to_H6M510_9_0 ),
    .H6M6(),
    .H6M7(\net_cnt_lcd_reg[7]_H6E7_to_H6M710_9_0 ),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(\net_cnt_lcd_reg[7]_H6E11_to_H6M1110_9_0 ),
    .H6W0(),
    .H6W1(\net_cnt_lcd_reg[4]_H6E1_to_H6W110_9_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(\net_Lut-U217_1_OUT6_to_OUT_E610_9_0 ),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(\net_Lut-U201_0_0_V6S0_to_V6M010_9_0 ),
    .V6M1(\net_Lut-U201_0_0_V6S1_to_V6M110_9_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(\net_cnt_lcd_reg[5]_V6S4_to_V6M410_9_0 ),
    .V6M5(),
    .V6M6(\net_cnt_lcd_reg[6]_V6S6_to_V6M610_9_0 ),
    .V6M7(),
    .V6M8(\net_Lut-U201_0_0_V6S8_to_V6M810_9_0 ),
    .V6M9(),
    .V6M10(\net_cnt_lcd_reg[5]_V6S10_to_V6M1010_9_0 ),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[7]_S0_F_B1_to_F110_9_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[6]_S0_F_B2_to_F210_9_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[0]_S0_F_B3_to_F310_9_0 ),
    .S0_F_B4(\net_Lut-U217_1_S0_F_B4_to_F410_9_0 ),
    .S0_G_B1(\net_cnt_lcd_reg[7]_S0_G_B1_to_G110_9_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[6]_S0_G_B2_to_G210_9_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[0]_S0_G_B3_to_G310_9_0 ),
    .S0_G_B4(\net_cnt_lcd_reg[5]_S0_G_B4_to_G410_9_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U152_0_0_X_to_S0_X10_9_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U170_0_Y_to_S0_Y10_9_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[5]_S1_F_B1_to_F110_9_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[3]_S1_F_B2_to_F210_9_0 ),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G110_9_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[3]_S1_G_B2_to_G210_9_0 ),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U227_0_X_to_S1_X10_9_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U161_0_0_Y_to_S1_Y10_9_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_10_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_h6w1.CONF = "0010";
  defparam GSB_CNT_10_10_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_h6w2.CONF = "0010";
  defparam GSB_CNT_10_10_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_10_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_10_0_inst.sps_n0.CONF = "01";
  defparam GSB_CNT_10_10_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n10.CONF = "10";
  defparam GSB_CNT_10_10_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_n6.CONF = "10";
  defparam GSB_CNT_10_10_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_n9.CONF = "10";
  defparam GSB_CNT_10_10_0_inst.sps_out0.CONF = "001011";
  defparam GSB_CNT_10_10_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_out2.CONF = "001011";
  defparam GSB_CNT_10_10_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_10_10_0_inst.sps_out4.CONF = "011101";
  defparam GSB_CNT_10_10_0_inst.sps_out5.CONF = "011101";
  defparam GSB_CNT_10_10_0_inst.sps_out6.CONF = "000111";
  defparam GSB_CNT_10_10_0_inst.sps_out7.CONF = "011110";
  defparam GSB_CNT_10_10_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s0_f_b1.CONF = "010101111";
  defparam GSB_CNT_10_10_0_inst.sps_s0_f_b2.CONF = "011111110";
  defparam GSB_CNT_10_10_0_inst.sps_s0_f_b3.CONF = "010110111";
  defparam GSB_CNT_10_10_0_inst.sps_s0_f_b4.CONF = "001111110";
  defparam GSB_CNT_10_10_0_inst.sps_s0_g_b1.CONF = "001000";
  defparam GSB_CNT_10_10_0_inst.sps_s0_g_b2.CONF = "001100";
  defparam GSB_CNT_10_10_0_inst.sps_s0_g_b3.CONF = "001111";
  defparam GSB_CNT_10_10_0_inst.sps_s0_g_b4.CONF = "010010";
  defparam GSB_CNT_10_10_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s17.CONF = "10";
  defparam GSB_CNT_10_10_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s1_f_b1.CONF = "010111101";
  defparam GSB_CNT_10_10_0_inst.sps_s1_f_b2.CONF = "011110111";
  defparam GSB_CNT_10_10_0_inst.sps_s1_f_b3.CONF = "011101111";
  defparam GSB_CNT_10_10_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_10_0_inst.sps_s1_g_b1.CONF = "011000";
  defparam GSB_CNT_10_10_0_inst.sps_s1_g_b2.CONF = "010010";
  defparam GSB_CNT_10_10_0_inst.sps_s1_g_b3.CONF = "010010";
  defparam GSB_CNT_10_10_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_10_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_v6n2.CONF = "0001";
  defparam GSB_CNT_10_10_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_10_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_10_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_w13.CONF = "0";
  defparam GSB_CNT_10_10_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w22.CONF = "10";
  defparam GSB_CNT_10_10_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_10_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e2_w2.CONF = "0";
  defparam GSB_CNT_10_10_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n11_w12.CONF = "0";
  defparam GSB_CNT_10_10_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n23_w0.CONF = "0";
  defparam GSB_CNT_10_10_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n7_w8.CONF = "0";
  defparam GSB_CNT_10_10_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s13_n13.CONF = "0";
  defparam GSB_CNT_10_10_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s21_e23.CONF = "0";
  defparam GSB_CNT_10_10_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s2_e20.CONF = "0";
  defparam GSB_CNT_10_10_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s9_e11.CONF = "0";
  defparam GSB_CNT_10_10_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_10_0_inst.switch_s9_w15.CONF = "0";
  GSB_CNT GSB_CNT_10_10_0_inst (
    .E0(),
    .E1(),
    .E2(\net_cnt_lcd_reg[4]_W2_to_E210_10_0 ),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(\net_cnt_lcd_reg[2]_W11_to_E1110_10_0 ),
    .E12(),
    .E13(),
    .E14(),
    .E15(\net_cnt_lcd_reg[7]_W15_to_E1510_10_0 ),
    .E16(\net_cnt_lcd_reg[3]_W16_to_E1610_10_0 ),
    .E17(),
    .E18(\net_cnt_lcd_reg[0]_W18_to_E1810_10_0 ),
    .E19(),
    .E20(\net_cnt_lcd_reg[0]_W20_to_E2010_10_0 ),
    .E21(),
    .E22(),
    .E23(\net_cnt_lcd_reg[3]_W23_to_E2310_10_0 ),
    .N0(\net_Lut-U224_0_0_N0_to_S09_10_0 ),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(\net_Lut-U224_0_0_N6_to_S69_10_0 ),
    .N7(\net_Lut-U227_0_N7_to_S79_10_0 ),
    .N8(\net_Lut-U223_0_S8_to_N810_10_0 ),
    .N9(\net_Lut-U225_0_N9_to_S99_10_0 ),
    .N10(\net_Lut-U205_0_0_N10_to_S109_10_0 ),
    .N11(),
    .N12(),
    .N13(\net_Lut-U216_0_N13_to_S139_10_0 ),
    .N14(),
    .N15(),
    .N16(),
    .N17(\net_Lut-U208_0_S17_to_N1710_10_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(\net_cnt_lcd_reg[5]_N23_to_S239_10_0 ),
    .W0(\net_cnt_lcd_reg[5]_E0_to_W010_10_0 ),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(\net_Lut-U227_0_E8_to_W810_10_0 ),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_cnt_lcd_reg[6]_E12_to_W1210_10_0 ),
    .W13(\net_Lut-U154_0_W13_to_E1310_9_0 ),
    .W14(\net_cnt_lcd_reg[7]_E14_to_W1410_10_0 ),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(\net_cnt_lcd_reg[5]_E21_to_W2110_10_0 ),
    .W22(\net_Lut-U195_0_W22_to_E2210_9_0 ),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(\net_Lut-U216_0_N13_to_S1310_10_0 ),
    .S14(),
    .S15(),
    .S16(),
    .S17(\net_Lut-U217_1_S17_to_N1711_10_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(\net_cnt_lcd_reg[3]_S21_to_N2111_10_0 ),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(\net_Lut-U205_0_0_H6E1_to_H6M110_10_0 ),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_Lut-U225_0_H6W1_to_H6M110_7_0 ),
    .H6W2(\net_Lut-U225_0_H6W2_to_H6M210_7_0 ),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(\net_Lut-U217_1_OUT6_to_OUT_E610_9_0 ),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(\net_Lut-U225_0_V6N2_to_V6M27_10_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(\net_Lut-U154_0_V6S8_to_V6M810_10_0 ),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[5]_S0_F_B1_to_F110_10_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[4]_S0_F_B2_to_F210_10_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[2]_S0_F_B3_to_F310_10_0 ),
    .S0_F_B4(\net_cnt_lcd_reg[3]_S0_F_B4_to_F410_10_0 ),
    .S0_G_B1(\net_cnt_lcd_reg[4]_S0_G_B1_to_G110_10_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[7]_S0_G_B2_to_G210_10_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[6]_S0_G_B3_to_G310_10_0 ),
    .S0_G_B4(\net_cnt_lcd_reg[0]_S0_G_B4_to_G410_10_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U217_1_X_to_S0_X10_10_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U224_0_0_Y_to_S0_Y10_10_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[7]_S1_F_B1_to_F110_10_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[6]_S1_F_B2_to_F210_10_0 ),
    .S1_F_B3(\net_cnt_lcd_reg[0]_S1_F_B3_to_F310_10_0 ),
    .S1_F_B4(),
    .S1_G_B1(\net_cnt_lcd_reg[2]_S1_G_B1_to_G110_10_0 ),
    .S1_G_B2(\net_Lut-U223_0_S1_G_B2_to_G210_10_0 ),
    .S1_G_B3(\net_Lut-U208_0_S1_G_B3_to_G310_10_0 ),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U225_0_X_to_S1_X10_10_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U195_0_Y_to_S1_Y10_10_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_9_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_e6.CONF = "10";
  defparam GSB_CNT_9_9_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_h6w2.CONF = "0010";
  defparam GSB_CNT_9_9_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_9_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_9_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_out2.CONF = "000111";
  defparam GSB_CNT_9_9_0_inst.sps_out3.CONF = "011110";
  defparam GSB_CNT_9_9_0_inst.sps_out4.CONF = "001011";
  defparam GSB_CNT_9_9_0_inst.sps_out5.CONF = "001011";
  defparam GSB_CNT_9_9_0_inst.sps_out6.CONF = "011101";
  defparam GSB_CNT_9_9_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s0_f_b1.CONF = "100110111";
  defparam GSB_CNT_9_9_0_inst.sps_s0_f_b2.CONF = "011111101";
  defparam GSB_CNT_9_9_0_inst.sps_s0_f_b3.CONF = "001111110";
  defparam GSB_CNT_9_9_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_9_0_inst.sps_s0_g_b1.CONF = "001011";
  defparam GSB_CNT_9_9_0_inst.sps_s0_g_b2.CONF = "011010";
  defparam GSB_CNT_9_9_0_inst.sps_s0_g_b3.CONF = "100101";
  defparam GSB_CNT_9_9_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s15.CONF = "10";
  defparam GSB_CNT_9_9_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s1_f_b1.CONF = "011110111";
  defparam GSB_CNT_9_9_0_inst.sps_s1_f_b2.CONF = "010101111";
  defparam GSB_CNT_9_9_0_inst.sps_s1_f_b3.CONF = "001111101";
  defparam GSB_CNT_9_9_0_inst.sps_s1_f_b4.CONF = "001111101";
  defparam GSB_CNT_9_9_0_inst.sps_s1_g_b1.CONF = "011000";
  defparam GSB_CNT_9_9_0_inst.sps_s1_g_b2.CONF = "011011";
  defparam GSB_CNT_9_9_0_inst.sps_s1_g_b3.CONF = "100000";
  defparam GSB_CNT_9_9_0_inst.sps_s1_g_b4.CONF = "001010";
  defparam GSB_CNT_9_9_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_9_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_v6n1.CONF = "0100";
  defparam GSB_CNT_9_9_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_9_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_9_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w11.CONF = "10";
  defparam GSB_CNT_9_9_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w17.CONF = "10";
  defparam GSB_CNT_9_9_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_9_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e5_w5.CONF = "0";
  defparam GSB_CNT_9_9_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_e9_w9.CONF = "0";
  defparam GSB_CNT_9_9_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_n9_w10.CONF = "0";
  defparam GSB_CNT_9_9_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_9_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_9_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(\net_cnt_lcd_reg[2]_E5_to_W59_10_0 ),
    .E6(),
    .E7(),
    .E8(\net_Lut-U205_0_0_W8_to_E89_9_0 ),
    .E9(\net_Lut-U224_0_1_W9_to_E99_9_0 ),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(\net_Lut-U204_0_1_S8_to_N89_9_0 ),
    .N9(\net_cnt_lcd_reg[4]_S9_to_N99_9_0 ),
    .N10(),
    .N11(),
    .N12(),
    .N13(\net_Lut-U176_0_1_S13_to_N139_9_0 ),
    .N14(),
    .N15(),
    .N16(),
    .N17(\net_cnt_lcd_reg[6]_S17_to_N179_9_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(\net_Lut-U229_0_S22_to_N229_9_0 ),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(\net_cnt_lcd_reg[2]_E5_to_W59_9_0 ),
    .W6(),
    .W7(),
    .W8(),
    .W9(\net_Lut-U224_0_1_W9_to_E99_8_0 ),
    .W10(),
    .W11(\net_Lut-U151_0_W11_to_E119_8_0 ),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(\net_Lut-U230_0_0_W17_to_E179_8_0 ),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(\net_cnt_lcd_reg[3]_E23_to_W239_9_0 ),
    .S0(),
    .S1(\net_Lut-U152_0_0_N1_to_S19_9_0 ),
    .S2(),
    .S3(),
    .S4(),
    .S5(\net_cnt_lcd_reg[5]_N5_to_S59_9_0 ),
    .S6(),
    .S7(),
    .S8(),
    .S9(\net_Lut-U227_0_N9_to_S99_9_0 ),
    .S10(),
    .S11(),
    .S12(),
    .S13(\net_Lut-U154_0_N13_to_S139_9_0 ),
    .S14(\net_cnt_lcd_reg[0]_N14_to_S149_9_0 ),
    .S15(\net_Lut-U230_0_0_S15_to_N1510_9_0 ),
    .S16(),
    .S17(\net_cnt_lcd_reg[7]_N17_to_S179_9_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(\net_Lut-U144_0_0_H6E1_to_H6M19_9_0 ),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(\net_Lut-U230_0_0_H6W2_to_H6M29_6_0 ),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(\net_Lut-U153_0_OUT6_to_OUT_E69_8_0 ),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(\net_Lut-U144_0_0_V6N1_to_V6M16_9_0 ),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U154_0_S0_F_B1_to_F19_9_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[4]_S0_F_B2_to_F29_9_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[3]_S0_F_B3_to_F39_9_0 ),
    .S0_F_B4(),
    .S0_G_B1(\net_cnt_lcd_reg[7]_S0_G_B1_to_G19_9_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[6]_S0_G_B2_to_G29_9_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[0]_S0_G_B3_to_G39_9_0 ),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U154_1_X_to_S0_X9_9_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U230_0_0_Y_to_S0_Y9_9_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U205_0_0_S1_F_B1_to_F19_9_0 ),
    .S1_F_B2(\net_Lut-U204_0_1_S1_F_B2_to_F29_9_0 ),
    .S1_F_B3(\net_Lut-U154_1_S1_F_B3_to_F39_9_0 ),
    .S1_F_B4(\net_cnt_lcd_reg[5]_S1_F_B4_to_F49_9_0 ),
    .S1_G_B1(\net_Lut-U227_0_S1_G_B1_to_G19_9_0 ),
    .S1_G_B2(\net_Lut-U176_0_1_S1_G_B2_to_G29_9_0 ),
    .S1_G_B3(\net_Lut-U152_0_0_S1_G_B3_to_G39_9_0 ),
    .S1_G_B4(\net_Lut-U229_0_S1_G_B4_to_G49_9_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U153_0_X_to_S1_X9_9_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U151_0_Y_to_S1_Y9_9_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_e0.CONF = "10";
  defparam GSB_CNT_10_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e10.CONF = "10";
  defparam GSB_CNT_10_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_e17.CONF = "10";
  defparam GSB_CNT_10_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_e21.CONF = "01";
  defparam GSB_CNT_10_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_h6e0.CONF = "0010";
  defparam GSB_CNT_10_6_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_h6e11.CONF = "010";
  defparam GSB_CNT_10_6_0_inst.sps_h6e2.CONF = "0010";
  defparam GSB_CNT_10_6_0_inst.sps_h6e3.CONF = "0011";
  defparam GSB_CNT_10_6_0_inst.sps_h6e5.CONF = "010";
  defparam GSB_CNT_10_6_0_inst.sps_h6e7.CONF = "010";
  defparam GSB_CNT_10_6_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_h6w2.CONF = "0100";
  defparam GSB_CNT_10_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_6_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n1.CONF = "10";
  defparam GSB_CNT_10_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_n9.CONF = "10";
  defparam GSB_CNT_10_6_0_inst.sps_out0.CONF = "000111";
  defparam GSB_CNT_10_6_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_out3.CONF = "001011";
  defparam GSB_CNT_10_6_0_inst.sps_out4.CONF = "011101";
  defparam GSB_CNT_10_6_0_inst.sps_out5.CONF = "011110";
  defparam GSB_CNT_10_6_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s0_f_b1.CONF = "001101111";
  defparam GSB_CNT_10_6_0_inst.sps_s0_f_b2.CONF = "100110111";
  defparam GSB_CNT_10_6_0_inst.sps_s0_f_b3.CONF = "010111011";
  defparam GSB_CNT_10_6_0_inst.sps_s0_f_b4.CONF = "011110111";
  defparam GSB_CNT_10_6_0_inst.sps_s0_g_b1.CONF = "001100";
  defparam GSB_CNT_10_6_0_inst.sps_s0_g_b2.CONF = "001100";
  defparam GSB_CNT_10_6_0_inst.sps_s0_g_b3.CONF = "100000";
  defparam GSB_CNT_10_6_0_inst.sps_s0_g_b4.CONF = "010000";
  defparam GSB_CNT_10_6_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s14.CONF = "01";
  defparam GSB_CNT_10_6_0_inst.sps_s15.CONF = "10";
  defparam GSB_CNT_10_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s1_f_b1.CONF = "001110111";
  defparam GSB_CNT_10_6_0_inst.sps_s1_f_b2.CONF = "010111110";
  defparam GSB_CNT_10_6_0_inst.sps_s1_f_b3.CONF = "100111110";
  defparam GSB_CNT_10_6_0_inst.sps_s1_f_b4.CONF = "100110111";
  defparam GSB_CNT_10_6_0_inst.sps_s1_g_b1.CONF = "100000";
  defparam GSB_CNT_10_6_0_inst.sps_s1_g_b2.CONF = "001111";
  defparam GSB_CNT_10_6_0_inst.sps_s1_g_b3.CONF = "011101";
  defparam GSB_CNT_10_6_0_inst.sps_s1_g_b4.CONF = "001011";
  defparam GSB_CNT_10_6_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s4.CONF = "01";
  defparam GSB_CNT_10_6_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_6_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_w2.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e12_w12.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e1_w1.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n0_e20.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n23_w0.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n4_e0.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s12_n12.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s23_w1.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s2_w0.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s5_n5.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s7_w9.CONF = "0";
  defparam GSB_CNT_10_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_6_0_inst (
    .E0(\net_cnt_lcd_reg[5]_E0_to_W010_7_0 ),
    .E1(\net_cnt_lcd_reg[2]_E1_to_W110_7_0 ),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(\net_cnt_lcd_reg[4]_E10_to_W1010_7_0 ),
    .E11(),
    .E12(\net_Lut-U232_0_0_E12_to_W1210_7_0 ),
    .E13(),
    .E14(),
    .E15(\net_Lut-U225_0_W15_to_E1510_6_0 ),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(\net_cnt_lcd_reg[7]_E21_to_W2110_7_0 ),
    .E22(),
    .E23(),
    .N0(\net_cnt_lcd_reg[2]_S0_to_N010_6_0 ),
    .N1(\net_Lut-U121_2_N1_to_S19_6_0 ),
    .N2(),
    .N3(),
    .N4(),
    .N5(\net_cnt_lcd_reg[4]_S5_to_N510_6_0 ),
    .N6(),
    .N7(\net_cnt_lcd_reg[4]_S7_to_N710_6_0 ),
    .N8(),
    .N9(\net_Lut-U117_0_N9_to_S99_6_0 ),
    .N10(),
    .N11(),
    .N12(\net_cnt_lcd_reg[3]_S12_to_N1210_6_0 ),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(\net_Lut-U230_0_0_S18_to_N1810_6_0 ),
    .N19(),
    .N20(),
    .N21(),
    .N22(\net_Lut-U122_0_0_S22_to_N2210_6_0 ),
    .N23(\net_cnt_lcd_reg[1]_N23_to_S239_6_0 ),
    .W0(\net_cnt_lcd_reg[1]_E0_to_W010_6_0 ),
    .W1(\net_cnt_lcd_reg[2]_E1_to_W110_6_0 ),
    .W2(\net_cnt_lcd_reg[5]_W2_to_E210_5_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(\net_cnt_lcd_reg[1]_E9_to_W910_6_0 ),
    .W10(),
    .W11(\net_Lut-U123_0_0_E11_to_W1110_6_0 ),
    .W12(\net_Lut-U232_0_0_E12_to_W1210_6_0 ),
    .W13(),
    .W14(),
    .W15(\net_cnt_lcd_reg[3]_E15_to_W1510_6_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(\net_Lut-U186_0_N0_to_S010_6_0 ),
    .S1(\net_Lut-U124_0_0_N1_to_S110_6_0 ),
    .S2(\net_cnt_lcd_reg[1]_S2_to_N211_6_0 ),
    .S3(),
    .S4(\net_cnt_lcd_reg[5]_S4_to_N411_6_0 ),
    .S5(),
    .S6(),
    .S7(\net_cnt_lcd_reg[1]_S7_to_N711_6_0 ),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(\net_cnt_lcd_reg[3]_S12_to_N1211_6_0 ),
    .S13(\net_Lut-U123_2_0_N13_to_S1310_6_0 ),
    .S14(\net_cnt_lcd_reg[4]_S14_to_N1411_6_0 ),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(\net_cnt_lcd_reg[5]_H6E0_to_H6M010_9_0 ),
    .H6E1(),
    .H6E2(\net_cnt_lcd_reg[6]_H6E2_to_H6M210_9_0 ),
    .H6E3(\net_cnt_lcd_reg[5]_H6E3_to_H6M310_9_0 ),
    .H6E4(),
    .H6E5(\net_cnt_lcd_reg[5]_H6E5_to_H6M510_9_0 ),
    .H6E6(),
    .H6E7(\net_cnt_lcd_reg[7]_H6E7_to_H6M710_9_0 ),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(\net_cnt_lcd_reg[7]_H6E11_to_H6M1110_9_0 ),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(\net_cnt_lcd_reg[4]_V6S2_to_V6N210_6_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(\net_cnt_lcd_reg[5]_V6S0_to_V6M010_6_0 ),
    .V6M1(),
    .V6M2(\net_cnt_lcd_reg[6]_V6S2_to_V6M210_6_0 ),
    .V6M3(\net_cnt_lcd_reg[5]_V6S3_to_V6M310_6_0 ),
    .V6M4(\net_cnt_lcd_reg[5]_V6S4_to_V6M410_6_0 ),
    .V6M5(),
    .V6M6(\net_cnt_lcd_reg[7]_V6S6_to_V6M610_6_0 ),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(\net_cnt_lcd_reg[7]_V6S10_to_V6M1010_6_0 ),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U122_0_0_S0_F_B1_to_F110_6_0 ),
    .S0_F_B2(\net_Lut-U230_0_0_S0_F_B2_to_F210_6_0 ),
    .S0_F_B3(\net_Lut-U123_1_S0_F_B3_to_F310_6_0 ),
    .S0_F_B4(\net_cnt_lcd_reg[4]_S0_F_B4_to_F410_6_0 ),
    .S0_G_B1(\net_cnt_lcd_reg[2]_S0_G_B1_to_G110_6_0 ),
    .S0_G_B2(\net_Lut-U225_0_S0_G_B2_to_G210_6_0 ),
    .S0_G_B3(\net_Lut-U186_0_S0_G_B3_to_G310_6_0 ),
    .S0_G_B4(\net_Lut-U118_0_0_S0_G_B4_to_G410_6_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U121_2_X_to_S0_X10_6_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U117_0_Y_to_S0_Y10_6_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U123_0_0_S1_F_B1_to_F110_6_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[5]_S1_F_B2_to_F210_6_0 ),
    .S1_F_B3(\net_Lut-U124_0_0_S1_F_B3_to_F310_6_0 ),
    .S1_F_B4(\net_Lut-U123_2_0_S1_F_B4_to_F410_6_0 ),
    .S1_G_B1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G110_6_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[3]_S1_G_B2_to_G210_6_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[2]_S1_G_B3_to_G310_6_0 ),
    .S1_G_B4(\net_cnt_lcd_reg[4]_S1_G_B4_to_G410_6_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U123_1_X_to_S1_X10_6_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U118_0_0_Y_to_S1_Y10_6_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e23.CONF = "01";
  defparam GSB_CNT_7_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_e5.CONF = "10";
  defparam GSB_CNT_7_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_h6e0.CONF = "0001";
  defparam GSB_CNT_7_5_0_inst.sps_h6e1.CONF = "0001";
  defparam GSB_CNT_7_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_h6e3.CONF = "0010";
  defparam GSB_CNT_7_5_0_inst.sps_h6e5.CONF = "001";
  defparam GSB_CNT_7_5_0_inst.sps_h6e7.CONF = "001";
  defparam GSB_CNT_7_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_5_0_inst.sps_h6w0.CONF = "0010";
  defparam GSB_CNT_7_5_0_inst.sps_h6w1.CONF = "0010";
  defparam GSB_CNT_7_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_5_0_inst.sps_h6w6.CONF = "000";
  defparam GSB_CNT_7_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n1.CONF = "10";
  defparam GSB_CNT_7_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_out0.CONF = "100111";
  defparam GSB_CNT_7_5_0_inst.sps_out1.CONF = "101011";
  defparam GSB_CNT_7_5_0_inst.sps_out2.CONF = "001011";
  defparam GSB_CNT_7_5_0_inst.sps_out3.CONF = "101011";
  defparam GSB_CNT_7_5_0_inst.sps_out4.CONF = "000111";
  defparam GSB_CNT_7_5_0_inst.sps_out5.CONF = "000111";
  defparam GSB_CNT_7_5_0_inst.sps_out6.CONF = "000111";
  defparam GSB_CNT_7_5_0_inst.sps_out7.CONF = "100111";
  defparam GSB_CNT_7_5_0_inst.sps_s0.CONF = "0";
  defparam GSB_CNT_7_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s0_f_b1.CONF = "001110111";
  defparam GSB_CNT_7_5_0_inst.sps_s0_f_b2.CONF = "011111011";
  defparam GSB_CNT_7_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_5_0_inst.sps_s0_g_b1.CONF = "011100";
  defparam GSB_CNT_7_5_0_inst.sps_s0_g_b2.CONF = "100101";
  defparam GSB_CNT_7_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s10.CONF = "10";
  defparam GSB_CNT_7_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s15.CONF = "10";
  defparam GSB_CNT_7_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s19.CONF = "0";
  defparam GSB_CNT_7_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s1_clk_b.CONF = "101011";
  defparam GSB_CNT_7_5_0_inst.sps_s1_f_b1.CONF = "011101111";
  defparam GSB_CNT_7_5_0_inst.sps_s1_f_b2.CONF = "010111011";
  defparam GSB_CNT_7_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_5_0_inst.sps_s1_g_b1.CONF = "100000";
  defparam GSB_CNT_7_5_0_inst.sps_s1_g_b2.CONF = "010101";
  defparam GSB_CNT_7_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_s1_sr_b.CONF = "111011";
  defparam GSB_CNT_7_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_s22.CONF = "10";
  defparam GSB_CNT_7_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_s8.CONF = "01";
  defparam GSB_CNT_7_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_v6s10.CONF = "001";
  defparam GSB_CNT_7_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_5_0_inst.sps_v6s4.CONF = "001";
  defparam GSB_CNT_7_5_0_inst.sps_v6s6.CONF = "001";
  defparam GSB_CNT_7_5_0_inst.sps_v6s8.CONF = "001";
  defparam GSB_CNT_7_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w22.CONF = "10";
  defparam GSB_CNT_7_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_5_0_inst.sps_w9.CONF = "10";
  defparam GSB_CNT_7_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n19_e19.CONF = "0";
  defparam GSB_CNT_7_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_5_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(\net_cnt_lcd_reg[1]_E5_to_W57_6_0 ),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(\net_cnt_lcd_reg[6]_W19_to_E197_5_0 ),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(\net_cnt_lcd_reg[1]_S0_to_N08_5_0 ),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(\net_cnt_lcd_reg[1]_S8_to_N88_5_0 ),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(net_U113_N14_to_S147_5_0),
    .S15(\net_Lut-U232_0_0_S15_to_N158_5_0 ),
    .S16(),
    .S17(),
    .S18(),
    .S19(\net_Lut-U232_0_0_S19_to_N198_5_0 ),
    .S20(),
    .S21(),
    .S22(\net_cnt_lcd_reg[0]_S22_to_N228_5_0 ),
    .S23(),
    .H6E0(\net_cnt_lcd_reg[1]_H6E0_to_H6M07_8_0 ),
    .H6E1(\net_cnt_lcd_reg[1]_H6E1_to_H6W17_11_0 ),
    .H6E2(),
    .H6E3(\net_cnt_lcd_reg[0]_H6E3_to_H6M37_8_0 ),
    .H6E4(),
    .H6E5(\net_cnt_lcd_reg[0]_H6E5_to_H6M57_8_0 ),
    .H6E6(),
    .H6E7(\net_Lut-U232_0_0_H6E7_to_H6M77_8_0 ),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(\net_cnt_lcd_reg[1]_H6W0_to_LEFT_H6M07_2_0 ),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_Lut-U232_0_0_H6W6_to_LEFT_H6M67_2_0 ),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBB1_to_GCLK17_3_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(\net_cnt_lcd_reg[1]_V6S4_to_V6M410_5_0 ),
    .V6S5(),
    .V6S6(\net_Lut-U232_0_0_V6S6_to_V6M610_5_0 ),
    .V6S7(),
    .V6S8(\net_cnt_lcd_reg[1]_V6S8_to_V6M810_5_0 ),
    .V6S9(),
    .V6S10(\net_cnt_lcd_reg[0]_V6S10_to_V6M1010_5_0 ),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(net_rst_nInvLut_V6N1_to_V6B17_5_0),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[6]_S0_F_B1_to_F17_5_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[0]_S0_F_B2_to_F27_5_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_cnt_lcd_reg[0]_S0_G_B1_to_G17_5_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G27_5_0 ),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U232_0_0_X_to_S0_X7_5_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U149_0_Y_to_S0_Y7_5_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[0]_S1_F_B1_to_F17_5_0 ),
    .S1_F_B2(net_U113_S1_F_B2_to_F27_5_0),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(\net_Lut-U149_0_S1_G_B1_to_G17_5_0 ),
    .S1_G_B2(net_U113_S1_G_B2_to_G27_5_0),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK7_5_0 ),
    .S1_SR_B(net_rst_nInvLut_S1_SR_B_to_SR7_5_0),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(\net_cnt_lcd_reg[0]_XQ_to_S1_XQ7_5_0 ),
    .S1_YQ(\net_cnt_lcd_reg[1]_YQ_to_S1_YQ7_5_0 ),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_e7.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n0_e20.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n14_w19.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n19_e19.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n22_e18.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s11_w13.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s15_n15.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s18_e12.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s22_n22.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s5_e7.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s8_n8.CONF = "0";
  defparam GSB_CNT_8_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_5_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(\net_cnt_lcd_reg[3]_E12_to_W128_6_0 ),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(\net_cnt_lcd_reg[0]_E18_to_W188_6_0 ),
    .E19(\net_Lut-U232_0_0_E19_to_W198_6_0 ),
    .E20(\net_cnt_lcd_reg[1]_E20_to_W208_6_0 ),
    .E21(),
    .E22(),
    .E23(),
    .N0(\net_cnt_lcd_reg[1]_S0_to_N08_5_0 ),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(\net_cnt_lcd_reg[1]_S8_to_N88_5_0 ),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(net_U113_N14_to_S147_5_0),
    .N15(\net_Lut-U232_0_0_S15_to_N158_5_0 ),
    .N16(),
    .N17(),
    .N18(),
    .N19(\net_Lut-U232_0_0_S19_to_N198_5_0 ),
    .N20(),
    .N21(),
    .N22(\net_cnt_lcd_reg[0]_S22_to_N228_5_0 ),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(net_U113_E13_to_W138_5_0),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(net_U113_E19_to_W198_5_0),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(\net_Buf-pad-rst_n_S5_to_N59_5_0 ),
    .S6(),
    .S7(),
    .S8(\net_cnt_lcd_reg[1]_S8_to_N89_5_0 ),
    .S9(),
    .S10(),
    .S11(net_U113_S11_to_N119_5_0),
    .S12(),
    .S13(),
    .S14(),
    .S15(\net_Lut-U232_0_0_S15_to_N159_5_0 ),
    .S16(),
    .S17(),
    .S18(\net_cnt_lcd_reg[3]_N18_to_S188_5_0 ),
    .S19(),
    .S20(),
    .S21(),
    .S22(\net_cnt_lcd_reg[0]_S22_to_N229_5_0 ),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_Buf-pad-rst_n_V6S1_to_V6M18_5_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_e15.CONF = "10";
  defparam GSB_CNT_9_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_e17.CONF = "10";
  defparam GSB_CNT_9_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_h6e1.CONF = "0001";
  defparam GSB_CNT_9_6_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_h6w8.CONF = "000";
  defparam GSB_CNT_9_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_6_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_n20.CONF = "10";
  defparam GSB_CNT_9_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_n9.CONF = "10";
  defparam GSB_CNT_9_6_0_inst.sps_out0.CONF = "011101";
  defparam GSB_CNT_9_6_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_out2.CONF = "000111";
  defparam GSB_CNT_9_6_0_inst.sps_out3.CONF = "001011";
  defparam GSB_CNT_9_6_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_out5.CONF = "001011";
  defparam GSB_CNT_9_6_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_out7.CONF = "011110";
  defparam GSB_CNT_9_6_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_s0_f_b1.CONF = "001110111";
  defparam GSB_CNT_9_6_0_inst.sps_s0_f_b2.CONF = "100111110";
  defparam GSB_CNT_9_6_0_inst.sps_s0_f_b3.CONF = "001110111";
  defparam GSB_CNT_9_6_0_inst.sps_s0_f_b4.CONF = "011111110";
  defparam GSB_CNT_9_6_0_inst.sps_s0_g_b1.CONF = "001010";
  defparam GSB_CNT_9_6_0_inst.sps_s0_g_b2.CONF = "010010";
  defparam GSB_CNT_9_6_0_inst.sps_s0_g_b3.CONF = "100000";
  defparam GSB_CNT_9_6_0_inst.sps_s0_g_b4.CONF = "010011";
  defparam GSB_CNT_9_6_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s18.CONF = "10";
  defparam GSB_CNT_9_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_s1_f_b1.CONF = "010110111";
  defparam GSB_CNT_9_6_0_inst.sps_s1_f_b2.CONF = "001110111";
  defparam GSB_CNT_9_6_0_inst.sps_s1_f_b3.CONF = "100110111";
  defparam GSB_CNT_9_6_0_inst.sps_s1_f_b4.CONF = "100111110";
  defparam GSB_CNT_9_6_0_inst.sps_s1_g_b1.CONF = "100100";
  defparam GSB_CNT_9_6_0_inst.sps_s1_g_b2.CONF = "100111";
  defparam GSB_CNT_9_6_0_inst.sps_s1_g_b3.CONF = "110111";
  defparam GSB_CNT_9_6_0_inst.sps_s1_g_b4.CONF = "110111";
  defparam GSB_CNT_9_6_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_s22.CONF = "10";
  defparam GSB_CNT_9_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_v6n7.CONF = "000";
  defparam GSB_CNT_9_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_6_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e2_w2.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n0_e20.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_n0_w5.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n19_e19.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n1_e1.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n5_e5.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n7_e7.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s0_w2.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s12_w14.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s23_e21.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s5_n5.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s7_n7.CONF = "0";
  defparam GSB_CNT_9_6_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_6_0_inst (
    .E0(),
    .E1(\net_cnt_lcd_reg[5]_E1_to_W19_7_0 ),
    .E2(\net_cnt_lcd_reg[2]_E2_to_W29_7_0 ),
    .E3(),
    .E4(),
    .E5(\net_cnt_lcd_reg[4]_E5_to_W59_7_0 ),
    .E6(),
    .E7(\net_cnt_lcd_reg[4]_E7_to_W79_7_0 ),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(\net_cnt_lcd_reg[3]_E15_to_W159_7_0 ),
    .E16(),
    .E17(\net_Lut-U144_0_0_E17_to_W179_7_0 ),
    .E18(),
    .E19(\net_Lut-U115_0_0_W19_to_E199_6_0 ),
    .E20(\net_cnt_lcd_reg[5]_E20_to_W209_7_0 ),
    .E21(\net_cnt_lcd_reg[1]_E21_to_W219_7_0 ),
    .E22(),
    .E23(),
    .N0(\net_cnt_lcd_reg[5]_S0_to_N09_6_0 ),
    .N1(\net_cnt_lcd_reg[5]_S1_to_N19_6_0 ),
    .N2(\net_cnt_lcd_reg[5]_S2_to_N29_6_0 ),
    .N3(\net_cnt_lcd_reg[1]_S3_to_N39_6_0 ),
    .N4(),
    .N5(\net_cnt_lcd_reg[4]_S5_to_N59_6_0 ),
    .N6(),
    .N7(\net_cnt_lcd_reg[4]_S7_to_N79_6_0 ),
    .N8(),
    .N9(\net_Lut-U144_0_0_N9_to_S98_6_0 ),
    .N10(),
    .N11(\net_Lut-U191_1_S11_to_N119_6_0 ),
    .N12(\net_cnt_lcd_reg[7]_S12_to_N129_6_0 ),
    .N13(),
    .N14(),
    .N15(),
    .N16(\net_cnt_lcd_reg[0]_S16_to_N169_6_0 ),
    .N17(),
    .N18(),
    .N19(),
    .N20(\net_cnt_lcd_reg[3]_N20_to_S208_6_0 ),
    .N21(),
    .N22(\net_cnt_lcd_reg[1]_S22_to_N229_6_0 ),
    .N23(),
    .W0(),
    .W1(),
    .W2(\net_cnt_lcd_reg[2]_E2_to_W29_6_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(\net_cnt_lcd_reg[3]_E14_to_W149_6_0 ),
    .W15(\net_Lut-U232_0_0_E15_to_W159_6_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(\net_cnt_lcd_reg[2]_S0_to_N010_6_0 ),
    .S1(\net_Lut-U121_2_N1_to_S19_6_0 ),
    .S2(),
    .S3(),
    .S4(),
    .S5(\net_cnt_lcd_reg[4]_S5_to_N510_6_0 ),
    .S6(),
    .S7(\net_cnt_lcd_reg[4]_S7_to_N710_6_0 ),
    .S8(),
    .S9(\net_Lut-U117_0_N9_to_S99_6_0 ),
    .S10(),
    .S11(),
    .S12(\net_cnt_lcd_reg[3]_S12_to_N1210_6_0 ),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(\net_Lut-U230_0_0_S18_to_N1810_6_0 ),
    .S19(),
    .S20(),
    .S21(),
    .S22(\net_Lut-U122_0_0_S22_to_N2210_6_0 ),
    .S23(\net_cnt_lcd_reg[1]_N23_to_S239_6_0 ),
    .H6E0(),
    .H6E1(\net_Lut-U144_0_0_H6E1_to_H6M19_9_0 ),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(\net_Lut-U230_0_0_H6W2_to_H6M29_6_0 ),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(\net_cnt_lcd_reg[3]_LEFT_H6B7_to_H6W79_6_0 ),
    .H6W8(\net_Lut-U115_1_H6W8_to_H6M89_3_0 ),
    .H6W9(),
    .H6W10(),
    .H6W11(\net_cnt_lcd_reg[3]_LEFT_H6B11_to_H6W119_6_0 ),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(\net_Lut-U166_0_OUT0_to_OUT_W09_7_0 ),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(\net_cnt_lcd_reg[2]_OUT0_to_OUT_W09_6_0 ),
    .OUT_W1(\net_cnt_lcd_reg[3]_OUT1_to_OUT_W19_6_0 ),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(\net_Lut-U144_0_0_V6N7_to_V6M76_6_0 ),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U115_0_0_S0_F_B1_to_F19_6_0 ),
    .S0_F_B2(\net_Lut-U121_2_S0_F_B2_to_F29_6_0 ),
    .S0_F_B3(\net_Lut-U191_1_S0_F_B3_to_F39_6_0 ),
    .S0_F_B4(\net_Lut-U117_0_S0_F_B4_to_F49_6_0 ),
    .S0_G_B1(\net_cnt_lcd_reg[1]_S0_G_B1_to_G19_6_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[0]_S0_G_B2_to_G29_6_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[2]_S0_G_B3_to_G39_6_0 ),
    .S0_G_B4(\net_cnt_lcd_reg[3]_S0_G_B4_to_G49_6_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U115_1_X_to_S0_X9_6_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U144_0_0_Y_to_S0_Y9_6_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[4]_S1_F_B1_to_F19_6_0 ),
    .S1_F_B2(\net_Lut-U232_0_0_S1_F_B2_to_F29_6_0 ),
    .S1_F_B3(\net_cnt_lcd_reg[7]_S1_F_B3_to_F39_6_0 ),
    .S1_F_B4(\net_cnt_lcd_reg[5]_S1_F_B4_to_F49_6_0 ),
    .S1_G_B1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G19_6_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[5]_S1_G_B2_to_G29_6_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[2]_S1_G_B3_to_G39_6_0 ),
    .S1_G_B4(\net_cnt_lcd_reg[3]_S1_G_B4_to_G49_6_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U166_0_X_to_S1_X9_6_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U122_0_0_Y_to_S1_Y9_6_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e2.CONF = "0010";
  defparam GSB_CNT_8_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6e9.CONF = "001";
  defparam GSB_CNT_8_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n14.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n21.CONF = "10";
  defparam GSB_CNT_8_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_n9.CONF = "10";
  defparam GSB_CNT_8_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_out2.CONF = "001011";
  defparam GSB_CNT_8_8_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_8_8_0_inst.sps_out4.CONF = "011110";
  defparam GSB_CNT_8_8_0_inst.sps_out5.CONF = "001011";
  defparam GSB_CNT_8_8_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_out7.CONF = "000111";
  defparam GSB_CNT_8_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_f_b1.CONF = "101111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_f_b2.CONF = "100111110";
  defparam GSB_CNT_8_8_0_inst.sps_s0_f_b3.CONF = "010111011";
  defparam GSB_CNT_8_8_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_g_b1.CONF = "110111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_g_b2.CONF = "001000";
  defparam GSB_CNT_8_8_0_inst.sps_s0_g_b3.CONF = "001000";
  defparam GSB_CNT_8_8_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s15.CONF = "10";
  defparam GSB_CNT_8_8_0_inst.sps_s16.CONF = "01";
  defparam GSB_CNT_8_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_f_b1.CONF = "010111101";
  defparam GSB_CNT_8_8_0_inst.sps_s1_f_b2.CONF = "011101111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_f_b3.CONF = "001111101";
  defparam GSB_CNT_8_8_0_inst.sps_s1_f_b4.CONF = "100111110";
  defparam GSB_CNT_8_8_0_inst.sps_s1_g_b1.CONF = "110111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_g_b2.CONF = "001111";
  defparam GSB_CNT_8_8_0_inst.sps_s1_g_b3.CONF = "001010";
  defparam GSB_CNT_8_8_0_inst.sps_s1_g_b4.CONF = "010010";
  defparam GSB_CNT_8_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e11_w11.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n17_e17.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n2_e22.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n4_e0.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n6_w11.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s11_n11.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s12_e10.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s17_e19.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s17_w23.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s1_w7.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s5_e7.CONF = "0";
  defparam GSB_CNT_8_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_8_0_inst (
    .E0(\net_cnt_lcd_reg[0]_E0_to_W08_9_0 ),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(\net_Lut-U202_0_0_W6_to_E68_8_0 ),
    .E7(\net_cnt_lcd_reg[2]_E7_to_W78_9_0 ),
    .E8(),
    .E9(),
    .E10(\net_cnt_lcd_reg[4]_W10_to_E108_8_0 ),
    .E11(\net_cnt_lcd_reg[1]_E11_to_W118_9_0 ),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(\net_Lut-U204_0_1_W17_to_E178_8_0 ),
    .E18(),
    .E19(\net_cnt_lcd_reg[3]_E19_to_W198_9_0 ),
    .E20(),
    .E21(),
    .E22(\net_cnt_lcd_reg[1]_E22_to_W228_9_0 ),
    .E23(),
    .N0(),
    .N1(),
    .N2(\net_cnt_lcd_reg[1]_S2_to_N28_8_0 ),
    .N3(),
    .N4(\net_cnt_lcd_reg[0]_S4_to_N48_8_0 ),
    .N5(),
    .N6(\net_cnt_lcd_reg[1]_S6_to_N68_8_0 ),
    .N7(),
    .N8(),
    .N9(\net_Lut-U189_2_N9_to_S97_8_0 ),
    .N10(),
    .N11(\net_Lut-U201_0_0_S11_to_N118_8_0 ),
    .N12(),
    .N13(),
    .N14(\net_Lut-U209_0_0_N14_to_S147_8_0 ),
    .N15(),
    .N16(\net_Lut-U232_0_0_S16_to_N168_8_0 ),
    .N17(\net_Lut-U204_0_1_N17_to_S177_8_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(\net_Lut-U178_0_N21_to_S217_8_0 ),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(\net_Lut-U190_0_1_E5_to_W58_8_0 ),
    .W6(),
    .W7(\net_cnt_lcd_reg[4]_E7_to_W78_8_0 ),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(\net_Lut-U225_0_E14_to_W148_8_0 ),
    .W15(\net_cnt_lcd_reg[7]_E15_to_W158_8_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(\net_Lut-U188_0_0_E21_to_W218_8_0 ),
    .W22(),
    .W23(\net_cnt_lcd_reg[3]_W23_to_E238_7_0 ),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(\net_cnt_lcd_reg[2]_N4_to_S48_8_0 ),
    .S5(\net_cnt_lcd_reg[2]_N5_to_S58_8_0 ),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(\net_Lut-U201_0_0_S11_to_N119_8_0 ),
    .S12(\net_cnt_lcd_reg[4]_S12_to_N129_8_0 ),
    .S13(),
    .S14(),
    .S15(),
    .S16(\net_Lut-U170_1_S16_to_N169_8_0 ),
    .S17(\net_cnt_lcd_reg[3]_N17_to_S178_8_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(\net_Lut-U209_0_0_H6E9_to_H6M98_11_0 ),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(\net_Lut-U213_0_0_OUT1_to_OUT_W18_8_0 ),
    .OUT_E6(\net_Lut-U180_0_0_OUT6_to_OUT_E68_8_0 ),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(\net_Lut-U170_1_V6N2_to_V6M28_8_0 ),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U189_2_S0_F_B1_to_F18_8_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[4]_S0_F_B2_to_F28_8_0 ),
    .S0_F_B3(\net_Lut-U179_2_S0_F_B3_to_F38_8_0 ),
    .S0_F_B4(),
    .S0_G_B1(\net_Lut-U213_0_0_S0_G_B1_to_G18_8_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[2]_S0_G_B2_to_G28_8_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[3]_S0_G_B3_to_G38_8_0 ),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U178_0_X_to_S0_X8_8_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U209_0_0_Y_to_S0_Y8_8_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U225_0_S1_F_B1_to_F18_8_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[2]_S1_F_B2_to_F28_8_0 ),
    .S1_F_B3(\net_Lut-U202_0_0_S1_F_B3_to_F38_8_0 ),
    .S1_F_B4(\net_Lut-U190_0_1_S1_F_B4_to_F48_8_0 ),
    .S1_G_B1(\net_Lut-U180_0_0_S1_G_B1_to_G18_8_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[7]_S1_G_B2_to_G28_8_0 ),
    .S1_G_B3(\net_Lut-U232_0_0_S1_G_B3_to_G38_8_0 ),
    .S1_G_B4(\net_Lut-U188_0_0_S1_G_B4_to_G48_8_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U189_2_X_to_S1_X8_8_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U179_2_Y_to_S1_Y8_8_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_11_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_h6e0.CONF = "0101";
  defparam GSB_CNT_7_11_0_inst.sps_h6e1.CONF = "0101";
  defparam GSB_CNT_7_11_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_11_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_11_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n19.CONF = "01";
  defparam GSB_CNT_7_11_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s4.CONF = "01";
  defparam GSB_CNT_7_11_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_s8.CONF = "01";
  defparam GSB_CNT_7_11_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_11_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_11_0_inst.sps_v6s3.CONF = "0010";
  defparam GSB_CNT_7_11_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_11_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w5.CONF = "01";
  defparam GSB_CNT_7_11_0_inst.sps_w6.CONF = "10";
  defparam GSB_CNT_7_11_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_11_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n19_w20.CONF = "0";
  defparam GSB_CNT_7_11_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_11_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_11_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(\net_cnt_lcd_reg[1]_W5_to_E57_10_0 ),
    .W6(\net_cnt_lcd_reg[1]_W6_to_E67_10_0 ),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(\net_cnt_lcd_reg[0]_W20_to_E207_10_0 ),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(\net_cnt_lcd_reg[1]_S4_to_N48_11_0 ),
    .S5(),
    .S6(),
    .S7(),
    .S8(\net_cnt_lcd_reg[1]_S8_to_N88_11_0 ),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(\net_cnt_lcd_reg[1]_H6E0_to_H6M07_8_0 ),
    .H6W1(\net_cnt_lcd_reg[1]_H6E1_to_H6W17_11_0 ),
    .H6W2(),
    .H6W3(\net_cnt_lcd_reg[0]_H6E3_to_H6M37_8_0 ),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(\net_cnt_lcd_reg[0]_V6S3_to_V6M310_11_0 ),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_11_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_h6e3.CONF = "0011";
  defparam GSB_CNT_10_11_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_11_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_11_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s6.CONF = "01";
  defparam GSB_CNT_10_11_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_11_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_11_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_11_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w18.CONF = "10";
  defparam GSB_CNT_10_11_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_w20.CONF = "01";
  defparam GSB_CNT_10_11_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_11_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e15_w15.CONF = "0";
  defparam GSB_CNT_10_11_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e2_w2.CONF = "0";
  defparam GSB_CNT_10_11_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n18_w23.CONF = "0";
  defparam GSB_CNT_10_11_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n6_w11.CONF = "0";
  defparam GSB_CNT_10_11_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s18_n18.CONF = "0";
  defparam GSB_CNT_10_11_0_inst.switch_s18_w16.CONF = "0";
  defparam GSB_CNT_10_11_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_11_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_11_0_inst (
    .E0(),
    .E1(),
    .E2(\net_cnt_lcd_reg[4]_W2_to_E210_11_0 ),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(\net_cnt_lcd_reg[7]_W15_to_E1510_11_0 ),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(\net_cnt_lcd_reg[2]_S6_to_N610_11_0 ),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(\net_cnt_lcd_reg[3]_S18_to_N1810_11_0 ),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(\net_cnt_lcd_reg[4]_W2_to_E210_10_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(\net_cnt_lcd_reg[2]_W11_to_E1110_10_0 ),
    .W12(),
    .W13(),
    .W14(),
    .W15(\net_cnt_lcd_reg[7]_W15_to_E1510_10_0 ),
    .W16(\net_cnt_lcd_reg[3]_W16_to_E1610_10_0 ),
    .W17(),
    .W18(\net_cnt_lcd_reg[0]_W18_to_E1810_10_0 ),
    .W19(),
    .W20(\net_cnt_lcd_reg[0]_W20_to_E2010_10_0 ),
    .W21(),
    .W22(),
    .W23(\net_cnt_lcd_reg[3]_W23_to_E2310_10_0 ),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(\net_cnt_lcd_reg[1]_S6_to_N611_11_0 ),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(\net_cnt_lcd_reg[1]_H6E5_to_H6M510_8_0 ),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(\net_cnt_lcd_reg[0]_V6S3_to_V6M310_11_0 ),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_e0.CONF = "10";
  defparam GSB_CNT_10_8_0_inst.sps_e1.CONF = "01";
  defparam GSB_CNT_10_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e19.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_e6.CONF = "10";
  defparam GSB_CNT_10_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_h6w10.CONF = "000";
  defparam GSB_CNT_10_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_h6w3.CONF = "0001";
  defparam GSB_CNT_10_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n5.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_out2.CONF = "001011";
  defparam GSB_CNT_10_8_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_out6.CONF = "011101";
  defparam GSB_CNT_10_8_0_inst.sps_out7.CONF = "011110";
  defparam GSB_CNT_10_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_s0_f_b1.CONF = "011111110";
  defparam GSB_CNT_10_8_0_inst.sps_s0_f_b2.CONF = "001111011";
  defparam GSB_CNT_10_8_0_inst.sps_s0_f_b3.CONF = "001101111";
  defparam GSB_CNT_10_8_0_inst.sps_s0_f_b4.CONF = "001111110";
  defparam GSB_CNT_10_8_0_inst.sps_s0_g_b1.CONF = "001101";
  defparam GSB_CNT_10_8_0_inst.sps_s0_g_b2.CONF = "010111";
  defparam GSB_CNT_10_8_0_inst.sps_s0_g_b3.CONF = "001010";
  defparam GSB_CNT_10_8_0_inst.sps_s0_g_b4.CONF = "001000";
  defparam GSB_CNT_10_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s16.CONF = "10";
  defparam GSB_CNT_10_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_s1_f_b1.CONF = "101111111";
  defparam GSB_CNT_10_8_0_inst.sps_s1_f_b2.CONF = "010111101";
  defparam GSB_CNT_10_8_0_inst.sps_s1_f_b3.CONF = "001111101";
  defparam GSB_CNT_10_8_0_inst.sps_s1_f_b4.CONF = "010111110";
  defparam GSB_CNT_10_8_0_inst.sps_s1_g_b1.CONF = "001101";
  defparam GSB_CNT_10_8_0_inst.sps_s1_g_b2.CONF = "100000";
  defparam GSB_CNT_10_8_0_inst.sps_s1_g_b3.CONF = "110111";
  defparam GSB_CNT_10_8_0_inst.sps_s1_g_b4.CONF = "110111";
  defparam GSB_CNT_10_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s4.CONF = "10";
  defparam GSB_CNT_10_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e13_w13.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e3_w3.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n16_e12.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.switch_n16_w21.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n19_w20.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_n9_e9.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s14_w12.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s4_w6.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.switch_s5_e7.CONF = "0";
  defparam GSB_CNT_10_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_8_0_inst (
    .E0(\net_cnt_lcd_reg[0]_E0_to_W010_9_0 ),
    .E1(\net_cnt_lcd_reg[1]_E1_to_W110_9_0 ),
    .E2(),
    .E3(\net_Lut-U201_0_0_W3_to_E310_8_0 ),
    .E4(),
    .E5(),
    .E6(),
    .E7(\net_Lut-U201_0_0_W7_to_E710_8_0 ),
    .E8(),
    .E9(\net_Lut-U161_0_0_W9_to_E910_8_0 ),
    .E10(\net_cnt_lcd_reg[4]_W10_to_E1010_8_0 ),
    .E11(),
    .E12(\net_cnt_lcd_reg[3]_E12_to_W1210_9_0 ),
    .E13(\net_Lut-U201_0_0_W13_to_E1310_8_0 ),
    .E14(),
    .E15(),
    .E16(\net_Lut-U230_0_0_W16_to_E1610_8_0 ),
    .E17(),
    .E18(),
    .E19(\net_cnt_lcd_reg[0]_E19_to_W1910_9_0 ),
    .E20(),
    .E21(),
    .E22(\net_Lut-U195_0_W22_to_E2210_8_0 ),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(\net_cnt_lcd_reg[1]_N5_to_S59_8_0 ),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(\net_Lut-U164_0_0_S12_to_N1210_8_0 ),
    .N13(),
    .N14(),
    .N15(),
    .N16(\net_cnt_lcd_reg[3]_S16_to_N1610_8_0 ),
    .N17(),
    .N18(),
    .N19(\net_Lut-U230_0_0_S19_to_N1910_8_0 ),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(\net_cnt_lcd_reg[5]_E0_to_W010_8_0 ),
    .W1(),
    .W2(),
    .W3(\net_Lut-U201_0_0_W3_to_E310_7_0 ),
    .W4(),
    .W5(),
    .W6(\net_cnt_lcd_reg[1]_W6_to_E610_7_0 ),
    .W7(\net_Lut-U205_0_0_E7_to_W710_8_0 ),
    .W8(\net_Lut-U159_0_0_E8_to_W810_8_0 ),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_Lut-U205_0_0_E12_to_W1210_8_0 ),
    .W13(\net_Lut-U201_0_0_W13_to_E1310_7_0 ),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(\net_Lut-U230_0_0_W20_to_E2010_7_0 ),
    .W21(\net_cnt_lcd_reg[3]_W21_to_E2110_7_0 ),
    .W22(),
    .W23(),
    .S0(\net_Lut-U196_4_N0_to_S010_8_0 ),
    .S1(),
    .S2(),
    .S3(),
    .S4(\net_cnt_lcd_reg[1]_S4_to_N411_8_0 ),
    .S5(\net_Lut-U201_0_0_S5_to_N511_8_0 ),
    .S6(),
    .S7(\net_Lut-U215_0_0_N7_to_S710_8_0 ),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(\net_Lut-U170_1_N12_to_S1210_8_0 ),
    .S13(),
    .S14(\net_Lut-U205_0_0_S14_to_N1411_8_0 ),
    .S15(),
    .S16(\net_Lut-U232_0_0_S16_to_N1611_8_0 ),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(\net_cnt_lcd_reg[1]_H6E5_to_H6M510_8_0 ),
    .H6M6(),
    .H6M7(\net_Lut-U232_0_0_H6E7_to_H6M710_8_0 ),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(\net_Lut-U195_1_H6W3_to_H6M310_5_0 ),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(\net_Lut-U157_1_H6W10_to_LEFT_H6E1010_2_0 ),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(\net_Lut-U196_6_1_OUT0_to_OUT_W010_8_0 ),
    .OUT_W1(\net_Lut-U196_7_1_OUT1_to_OUT_W110_8_0 ),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(\net_cnt_lcd_reg[1]_V6S0_to_V6M010_8_0 ),
    .V6M1(),
    .V6M2(),
    .V6M3(\net_cnt_lcd_reg[0]_V6S3_to_V6M310_8_0 ),
    .V6M4(\net_cnt_lcd_reg[0]_V6S4_to_V6M410_8_0 ),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U161_0_0_S0_F_B1_to_F110_8_0 ),
    .S0_F_B2(\net_Lut-U215_0_0_S0_F_B2_to_F210_8_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[4]_S0_F_B3_to_F310_8_0 ),
    .S0_F_B4(\net_Lut-U230_0_0_S0_F_B4_to_F410_8_0 ),
    .S0_G_B1(\net_Lut-U205_0_0_S0_G_B1_to_G110_8_0 ),
    .S0_G_B2(\net_Lut-U164_0_0_S0_G_B2_to_G210_8_0 ),
    .S0_G_B3(\net_Lut-U159_0_0_S0_G_B3_to_G310_8_0 ),
    .S0_G_B4(\net_Lut-U230_0_0_S0_G_B4_to_G410_8_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U160_0_X_to_S0_X10_8_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U158_0_Y_to_S0_Y10_8_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U160_0_S1_F_B1_to_F110_8_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[5]_S1_F_B2_to_F210_8_0 ),
    .S1_F_B3(\net_Lut-U158_0_S1_F_B3_to_F310_8_0 ),
    .S1_F_B4(\net_Lut-U170_1_S1_F_B4_to_F410_8_0 ),
    .S1_G_B1(\net_Lut-U195_0_S1_G_B1_to_G110_8_0 ),
    .S1_G_B2(\net_Lut-U196_4_S1_G_B2_to_G210_8_0 ),
    .S1_G_B3(\net_Lut-U196_6_1_S1_G_B3_to_G310_8_0 ),
    .S1_G_B4(\net_Lut-U196_7_1_S1_G_B4_to_G410_8_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U157_1_X_to_S1_X10_8_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U195_1_Y_to_S1_Y10_8_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e14.CONF = "0";
  defparam GSB_CNT_9_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_e2.CONF = "0";
  defparam GSB_CNT_9_5_0_inst.sps_e20.CONF = "0";
  defparam GSB_CNT_9_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_h6e0.CONF = "0011";
  defparam GSB_CNT_9_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_h6e11.CONF = "001";
  defparam GSB_CNT_9_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_h6e5.CONF = "001";
  defparam GSB_CNT_9_5_0_inst.sps_h6e7.CONF = "001";
  defparam GSB_CNT_9_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_h6w10.CONF = "000";
  defparam GSB_CNT_9_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_5_0_inst.sps_h6w6.CONF = "000";
  defparam GSB_CNT_9_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_5_0_inst.sps_n0.CONF = "01";
  defparam GSB_CNT_9_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_n18.CONF = "10";
  defparam GSB_CNT_9_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_out0.CONF = "001101";
  defparam GSB_CNT_9_5_0_inst.sps_out1.CONF = "001110";
  defparam GSB_CNT_9_5_0_inst.sps_out2.CONF = "011101";
  defparam GSB_CNT_9_5_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_9_5_0_inst.sps_out4.CONF = "001110";
  defparam GSB_CNT_9_5_0_inst.sps_out5.CONF = "011101";
  defparam GSB_CNT_9_5_0_inst.sps_out6.CONF = "001110";
  defparam GSB_CNT_9_5_0_inst.sps_out7.CONF = "011110";
  defparam GSB_CNT_9_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_9_5_0_inst.sps_s0_f_b1.CONF = "001011111";
  defparam GSB_CNT_9_5_0_inst.sps_s0_f_b2.CONF = "010111011";
  defparam GSB_CNT_9_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_5_0_inst.sps_s0_g_b1.CONF = "100111";
  defparam GSB_CNT_9_5_0_inst.sps_s0_g_b2.CONF = "010101";
  defparam GSB_CNT_9_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s0_sr_b.CONF = "001101";
  defparam GSB_CNT_9_5_0_inst.sps_s1.CONF = "10";
  defparam GSB_CNT_9_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s14.CONF = "10";
  defparam GSB_CNT_9_5_0_inst.sps_s15.CONF = "10";
  defparam GSB_CNT_9_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s17.CONF = "10";
  defparam GSB_CNT_9_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s1_f_b1.CONF = "100111011";
  defparam GSB_CNT_9_5_0_inst.sps_s1_f_b2.CONF = "011110111";
  defparam GSB_CNT_9_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_5_0_inst.sps_s1_g_b1.CONF = "011100";
  defparam GSB_CNT_9_5_0_inst.sps_s1_g_b2.CONF = "010010";
  defparam GSB_CNT_9_5_0_inst.sps_s1_g_b3.CONF = "011100";
  defparam GSB_CNT_9_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_s3.CONF = "10";
  defparam GSB_CNT_9_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_v6n0.CONF = "0001";
  defparam GSB_CNT_9_5_0_inst.sps_v6n1.CONF = "0001";
  defparam GSB_CNT_9_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_5_0_inst.sps_v6n2.CONF = "0001";
  defparam GSB_CNT_9_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_v6n5.CONF = "000";
  defparam GSB_CNT_9_5_0_inst.sps_v6n7.CONF = "000";
  defparam GSB_CNT_9_5_0_inst.sps_v6n9.CONF = "000";
  defparam GSB_CNT_9_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_5_0_inst.sps_v6s2.CONF = "0000";
  defparam GSB_CNT_9_5_0_inst.sps_v6s3.CONF = "0000";
  defparam GSB_CNT_9_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_w10.CONF = "10";
  defparam GSB_CNT_9_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n15_e15.CONF = "0";
  defparam GSB_CNT_9_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n22_e18.CONF = "0";
  defparam GSB_CNT_9_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s14_w12.CONF = "0";
  defparam GSB_CNT_9_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s22_w20.CONF = "0";
  defparam GSB_CNT_9_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_5_0_inst (
    .E0(),
    .E1(),
    .E2(\net_cnt_lcd_reg[2]_E2_to_W29_6_0 ),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(\net_cnt_lcd_reg[3]_E14_to_W149_6_0 ),
    .E15(\net_Lut-U232_0_0_E15_to_W159_6_0 ),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(\net_Buf-pad-rst_n_S5_to_N59_5_0 ),
    .N6(),
    .N7(),
    .N8(\net_cnt_lcd_reg[1]_S8_to_N89_5_0 ),
    .N9(),
    .N10(),
    .N11(net_U113_S11_to_N119_5_0),
    .N12(),
    .N13(),
    .N14(),
    .N15(\net_Lut-U232_0_0_S15_to_N159_5_0 ),
    .N16(),
    .N17(),
    .N18(\net_cnt_lcd_reg[3]_N18_to_S188_5_0 ),
    .N19(),
    .N20(),
    .N21(),
    .N22(\net_cnt_lcd_reg[0]_S22_to_N229_5_0 ),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(net_rst_nInvLut_W10_to_E109_4_0),
    .W11(),
    .W12(\net_Lut-U162_1_W12_to_E129_4_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(\net_Lut-U195_1_W20_to_E209_4_0 ),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(\net_cnt_lcd_reg[2]_S1_to_N110_5_0 ),
    .S2(),
    .S3(\net_cnt_lcd_reg[2]_S3_to_N310_5_0 ),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(\net_Lut-U145_0_N13_to_S139_5_0 ),
    .S14(),
    .S15(\net_cnt_lcd_reg[3]_S15_to_N1510_5_0 ),
    .S16(),
    .S17(\net_cnt_lcd_reg[3]_S17_to_N1710_5_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(\net_Lut-U195_1_N22_to_S229_5_0 ),
    .S23(net_U113_N23_to_S239_5_0),
    .H6E0(\net_cnt_lcd_reg[2]_H6E0_to_H6M09_8_0 ),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(\net_cnt_lcd_reg[2]_H6E5_to_H6M59_8_0 ),
    .H6E6(),
    .H6E7(\net_cnt_lcd_reg[3]_H6E7_to_H6M79_8_0 ),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(\net_cnt_lcd_reg[3]_H6E11_to_H6M119_8_0 ),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(\net_Lut-U162_1_H6W6_to_H6M69_5_0 ),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_cnt_lcd_reg[3]_H6W6_to_LEFT_H6M69_2_0 ),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(\net_cnt_lcd_reg[3]_H6W10_to_LEFT_H6M109_2_0 ),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBD1_to_GCLK19_3_0 ),
    .GCLK0(),
    .OUT0(\net_cnt_lcd_reg[2]_OUT0_to_OUT_W09_6_0 ),
    .OUT1(\net_cnt_lcd_reg[3]_OUT1_to_OUT_W19_6_0 ),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(\net_cnt_lcd_reg[2]_V6N0_to_V6M06_5_0 ),
    .V6N1(net_rst_nInvLut_V6N1_to_V6B17_5_0),
    .V6N2(\net_cnt_lcd_reg[3]_V6N2_to_V6M26_5_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(\net_cnt_lcd_reg[3]_V6N5_to_V6M56_5_0 ),
    .V6N6(),
    .V6N7(net_rst_nInvLut_V6N7_to_V6M76_5_0),
    .V6N8(),
    .V6N9(net_rst_nInvLut_V6N9_to_V6M96_5_0),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(\net_cnt_lcd_reg[3]_V6S2_to_V6M212_5_0 ),
    .V6S3(\net_cnt_lcd_reg[3]_V6S3_to_V6M312_5_0 ),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U147_0_S0_F_B1_to_F19_5_0 ),
    .S0_F_B2(net_U113_S0_F_B2_to_F29_5_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Lut-U145_0_S0_G_B1_to_G19_5_0 ),
    .S0_G_B2(net_U113_S0_G_B2_to_G29_5_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK9_5_0 ),
    .S0_SR_B(net_rst_nInvLut_S0_SR_B_to_SR9_5_0),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_cnt_lcd_reg[2]_XQ_to_S0_XQ9_5_0 ),
    .S0_YQ(\net_cnt_lcd_reg[3]_YQ_to_S0_YQ9_5_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Buf-pad-rst_n_S1_F_B1_to_F19_5_0 ),
    .S1_F_B2(net_U113_S1_F_B2_to_F29_5_0),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(\net_cnt_lcd_reg[2]_S1_G_B1_to_G19_5_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[1]_S1_G_B2_to_G29_5_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[0]_S1_G_B3_to_G39_5_0 ),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(net_rst_nInvLut_X_to_S1_X9_5_0),
    .S1_XB(),
    .S1_Y(\net_Lut-U147_0_Y_to_S1_Y9_5_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_e0.CONF = "10";
  defparam GSB_CNT_10_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e11.CONF = "01";
  defparam GSB_CNT_10_5_0_inst.sps_e12.CONF = "10";
  defparam GSB_CNT_10_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_e21.CONF = "01";
  defparam GSB_CNT_10_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_e9.CONF = "01";
  defparam GSB_CNT_10_5_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_h6e5.CONF = "010";
  defparam GSB_CNT_10_5_0_inst.sps_h6e7.CONF = "010";
  defparam GSB_CNT_10_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n13.CONF = "10";
  defparam GSB_CNT_10_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n22.CONF = "10";
  defparam GSB_CNT_10_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_out3.CONF = "000111";
  defparam GSB_CNT_10_5_0_inst.sps_out4.CONF = "001011";
  defparam GSB_CNT_10_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s0_f_b1.CONF = "001111110";
  defparam GSB_CNT_10_5_0_inst.sps_s0_f_b2.CONF = "011101111";
  defparam GSB_CNT_10_5_0_inst.sps_s0_f_b3.CONF = "011110111";
  defparam GSB_CNT_10_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_5_0_inst.sps_s0_g_b1.CONF = "011111";
  defparam GSB_CNT_10_5_0_inst.sps_s0_g_b2.CONF = "011000";
  defparam GSB_CNT_10_5_0_inst.sps_s0_g_b3.CONF = "100011";
  defparam GSB_CNT_10_5_0_inst.sps_s0_g_b4.CONF = "001010";
  defparam GSB_CNT_10_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_w2.CONF = "0";
  defparam GSB_CNT_10_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n15_e15.CONF = "0";
  defparam GSB_CNT_10_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n1_e1.CONF = "0";
  defparam GSB_CNT_10_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n23_w0.CONF = "0";
  defparam GSB_CNT_10_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n3_w4.CONF = "0";
  defparam GSB_CNT_10_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s1_n1.CONF = "0";
  defparam GSB_CNT_10_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_5_0_inst (
    .E0(\net_cnt_lcd_reg[1]_E0_to_W010_6_0 ),
    .E1(\net_cnt_lcd_reg[2]_E1_to_W110_6_0 ),
    .E2(\net_cnt_lcd_reg[5]_W2_to_E210_5_0 ),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(\net_cnt_lcd_reg[1]_E9_to_W910_6_0 ),
    .E10(),
    .E11(\net_Lut-U123_0_0_E11_to_W1110_6_0 ),
    .E12(\net_Lut-U232_0_0_E12_to_W1210_6_0 ),
    .E13(),
    .E14(),
    .E15(\net_cnt_lcd_reg[3]_E15_to_W1510_6_0 ),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(\net_cnt_lcd_reg[2]_S1_to_N110_5_0 ),
    .N2(),
    .N3(\net_cnt_lcd_reg[2]_S3_to_N310_5_0 ),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(\net_Lut-U145_0_N13_to_S139_5_0 ),
    .N14(),
    .N15(\net_cnt_lcd_reg[3]_S15_to_N1510_5_0 ),
    .N16(),
    .N17(\net_cnt_lcd_reg[3]_S17_to_N1710_5_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(\net_Lut-U195_1_N22_to_S229_5_0 ),
    .N23(net_U113_N23_to_S239_5_0),
    .W0(net_U113_E0_to_W010_5_0),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(\net_cnt_lcd_reg[2]_S1_to_N111_5_0 ),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(\net_cnt_lcd_reg[1]_H6E5_to_H6M510_8_0 ),
    .H6E6(),
    .H6E7(\net_Lut-U232_0_0_H6E7_to_H6M710_8_0 ),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(\net_Lut-U195_1_H6W3_to_H6M310_5_0 ),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(\net_cnt_lcd_reg[1]_V6S4_to_V6M410_5_0 ),
    .V6M5(),
    .V6M6(\net_Lut-U232_0_0_V6S6_to_V6M610_5_0 ),
    .V6M7(),
    .V6M8(\net_cnt_lcd_reg[1]_V6S8_to_V6M810_5_0 ),
    .V6M9(),
    .V6M10(\net_cnt_lcd_reg[0]_V6S10_to_V6M1010_5_0 ),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[5]_S0_F_B1_to_F110_5_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[3]_S0_F_B2_to_F210_5_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[2]_S0_F_B3_to_F310_5_0 ),
    .S0_F_B4(),
    .S0_G_B1(\net_cnt_lcd_reg[3]_S0_G_B1_to_G110_5_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G210_5_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[0]_S0_G_B3_to_G310_5_0 ),
    .S0_G_B4(\net_cnt_lcd_reg[2]_S0_G_B4_to_G410_5_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U123_0_0_X_to_S0_X10_5_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U145_0_Y_to_S0_Y10_5_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_8_0_inst.sps_n0.CONF = "01";
  defparam GSB_CNT_11_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n12.CONF = "01";
  defparam GSB_CNT_11_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_out0.CONF = "011110";
  defparam GSB_CNT_11_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_out3.CONF = "001011";
  defparam GSB_CNT_11_8_0_inst.sps_out4.CONF = "011101";
  defparam GSB_CNT_11_8_0_inst.sps_out5.CONF = "000111";
  defparam GSB_CNT_11_8_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_f_b1.CONF = "100111011";
  defparam GSB_CNT_11_8_0_inst.sps_s0_f_b2.CONF = "100011111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_f_b3.CONF = "110111111";
  defparam GSB_CNT_11_8_0_inst.sps_s0_f_b4.CONF = "001111011";
  defparam GSB_CNT_11_8_0_inst.sps_s0_g_b1.CONF = "100101";
  defparam GSB_CNT_11_8_0_inst.sps_s0_g_b2.CONF = "100100";
  defparam GSB_CNT_11_8_0_inst.sps_s0_g_b3.CONF = "010000";
  defparam GSB_CNT_11_8_0_inst.sps_s0_g_b4.CONF = "011101";
  defparam GSB_CNT_11_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_f_b1.CONF = "010111110";
  defparam GSB_CNT_11_8_0_inst.sps_s1_f_b2.CONF = "001011111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_f_b3.CONF = "100111110";
  defparam GSB_CNT_11_8_0_inst.sps_s1_f_b4.CONF = "100110111";
  defparam GSB_CNT_11_8_0_inst.sps_s1_g_b1.CONF = "010011";
  defparam GSB_CNT_11_8_0_inst.sps_s1_g_b2.CONF = "001010";
  defparam GSB_CNT_11_8_0_inst.sps_s1_g_b3.CONF = "011101";
  defparam GSB_CNT_11_8_0_inst.sps_s1_g_b4.CONF = "011000";
  defparam GSB_CNT_11_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n2.CONF = "0001";
  defparam GSB_CNT_11_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w11.CONF = "10";
  defparam GSB_CNT_11_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w16.CONF = "10";
  defparam GSB_CNT_11_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e1_w1.CONF = "0";
  defparam GSB_CNT_11_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n16_e12.CONF = "0";
  defparam GSB_CNT_11_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n4_e0.CONF = "0";
  defparam GSB_CNT_11_8_0_inst.switch_n4_w9.CONF = "0";
  defparam GSB_CNT_11_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n7_e7.CONF = "0";
  defparam GSB_CNT_11_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_n9_e9.CONF = "0";
  defparam GSB_CNT_11_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s23_e21.CONF = "0";
  defparam GSB_CNT_11_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s4_e2.CONF = "0";
  defparam GSB_CNT_11_8_0_inst.switch_s4_n4.CONF = "0";
  defparam GSB_CNT_11_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_8_0_inst (
    .E0(\net_cnt_lcd_reg[1]_E0_to_W011_9_0 ),
    .E1(\net_Lut-U204_0_1_W1_to_E111_8_0 ),
    .E2(\net_cnt_lcd_reg[1]_E2_to_W211_9_0 ),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(\net_Lut-U215_0_0_W7_to_E711_8_0 ),
    .E8(),
    .E9(\net_Lut-U196_5_1_W9_to_E911_8_0 ),
    .E10(\net_cnt_lcd_reg[4]_W10_to_E1011_8_0 ),
    .E11(),
    .E12(\net_Lut-U232_0_0_E12_to_W1211_9_0 ),
    .E13(\net_Lut-U204_0_1_W13_to_E1311_8_0 ),
    .E14(),
    .E15(),
    .E16(),
    .E17(\net_Lut-U170_0_W17_to_E1711_8_0 ),
    .E18(),
    .E19(),
    .E20(),
    .E21(\net_Lut-U196_4_1_W21_to_E2111_8_0 ),
    .E22(\net_cnt_lcd_reg[5]_W22_to_E2211_8_0 ),
    .E23(),
    .N0(\net_Lut-U196_4_N0_to_S010_8_0 ),
    .N1(),
    .N2(),
    .N3(),
    .N4(\net_cnt_lcd_reg[1]_S4_to_N411_8_0 ),
    .N5(\net_Lut-U201_0_0_S5_to_N511_8_0 ),
    .N6(),
    .N7(\net_Lut-U215_0_0_N7_to_S710_8_0 ),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(\net_Lut-U170_1_N12_to_S1210_8_0 ),
    .N13(),
    .N14(\net_Lut-U205_0_0_S14_to_N1411_8_0 ),
    .N15(),
    .N16(\net_Lut-U232_0_0_S16_to_N1611_8_0 ),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(\net_Lut-U204_0_1_W1_to_E111_7_0 ),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(\net_Lut-U196_3_1_E6_to_W611_8_0 ),
    .W7(),
    .W8(),
    .W9(\net_cnt_lcd_reg[1]_W9_to_E911_7_0 ),
    .W10(),
    .W11(\net_Lut-U196_1_0_W11_to_E1111_7_0 ),
    .W12(),
    .W13(),
    .W14(\net_Lut-U196_1_E14_to_W1411_8_0 ),
    .W15(),
    .W16(\net_Lut-U196_0_1_W16_to_E1611_7_0 ),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(\net_cnt_lcd_reg[2]_N1_to_S111_8_0 ),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(\net_cnt_lcd_reg[3]_N13_to_S1311_8_0 ),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(\net_Lut-U202_0_0_OUT7_to_OUT_E711_8_0 ),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(\net_Lut-U170_1_V6N2_to_V6M28_8_0 ),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U205_0_0_S0_F_B1_to_F111_8_0 ),
    .S0_F_B2(\net_Lut-U204_0_1_S0_F_B2_to_F211_8_0 ),
    .S0_F_B3(\net_Lut-U202_0_0_S0_F_B3_to_F311_8_0 ),
    .S0_F_B4(\net_Lut-U201_0_0_S0_F_B4_to_F411_8_0 ),
    .S0_G_B1(\net_Lut-U205_0_0_S0_G_B1_to_G111_8_0 ),
    .S0_G_B2(\net_Lut-U204_0_1_S0_G_B2_to_G211_8_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[1]_S0_G_B3_to_G311_8_0 ),
    .S0_G_B4(\net_cnt_lcd_reg[5]_S0_G_B4_to_G411_8_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U196_0_1_X_to_S0_X11_8_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U196_1_0_Y_to_S0_Y11_8_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U170_0_S1_F_B1_to_F111_8_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[4]_S1_F_B2_to_F211_8_0 ),
    .S1_F_B3(\net_cnt_lcd_reg[2]_S1_F_B3_to_F311_8_0 ),
    .S1_F_B4(\net_cnt_lcd_reg[3]_S1_F_B4_to_F411_8_0 ),
    .S1_G_B1(\net_Lut-U196_1_S1_G_B1_to_G111_8_0 ),
    .S1_G_B2(\net_Lut-U196_3_1_S1_G_B2_to_G211_8_0 ),
    .S1_G_B3(\net_Lut-U196_4_1_S1_G_B3_to_G311_8_0 ),
    .S1_G_B4(\net_Lut-U196_5_1_S1_G_B4_to_G411_8_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U170_1_X_to_S1_X11_8_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U196_4_Y_to_S1_Y11_8_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_7_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e14.CONF = "0";
  defparam GSB_CNT_11_7_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_e6.CONF = "10";
  defparam GSB_CNT_11_7_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_7_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_7_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_out2.CONF = "001011";
  defparam GSB_CNT_11_7_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_11_7_0_inst.sps_out4.CONF = "000111";
  defparam GSB_CNT_11_7_0_inst.sps_out5.CONF = "011110";
  defparam GSB_CNT_11_7_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s0_f_b1.CONF = "100011111";
  defparam GSB_CNT_11_7_0_inst.sps_s0_f_b2.CONF = "001111101";
  defparam GSB_CNT_11_7_0_inst.sps_s0_f_b3.CONF = "011111101";
  defparam GSB_CNT_11_7_0_inst.sps_s0_f_b4.CONF = "001110111";
  defparam GSB_CNT_11_7_0_inst.sps_s0_g_b1.CONF = "010000";
  defparam GSB_CNT_11_7_0_inst.sps_s0_g_b2.CONF = "011011";
  defparam GSB_CNT_11_7_0_inst.sps_s0_g_b3.CONF = "001010";
  defparam GSB_CNT_11_7_0_inst.sps_s0_g_b4.CONF = "100000";
  defparam GSB_CNT_11_7_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_s12.CONF = "0";
  defparam GSB_CNT_11_7_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s1_f_b1.CONF = "010111011";
  defparam GSB_CNT_11_7_0_inst.sps_s1_f_b2.CONF = "100111011";
  defparam GSB_CNT_11_7_0_inst.sps_s1_f_b3.CONF = "011111101";
  defparam GSB_CNT_11_7_0_inst.sps_s1_f_b4.CONF = "010110111";
  defparam GSB_CNT_11_7_0_inst.sps_s1_g_b1.CONF = "100101";
  defparam GSB_CNT_11_7_0_inst.sps_s1_g_b2.CONF = "100101";
  defparam GSB_CNT_11_7_0_inst.sps_s1_g_b3.CONF = "011011";
  defparam GSB_CNT_11_7_0_inst.sps_s1_g_b4.CONF = "010111";
  defparam GSB_CNT_11_7_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_7_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_v6n2.CONF = "0100";
  defparam GSB_CNT_11_7_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_v6n5.CONF = "011";
  defparam GSB_CNT_11_7_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_7_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_7_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w11.CONF = "10";
  defparam GSB_CNT_11_7_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_7_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_e9_w9.CONF = "0";
  defparam GSB_CNT_11_7_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n20_e16.CONF = "0";
  defparam GSB_CNT_11_7_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_7_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_7_0_inst (
    .E0(),
    .E1(\net_Lut-U204_0_1_W1_to_E111_7_0 ),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(\net_Lut-U196_3_1_E6_to_W611_8_0 ),
    .E7(),
    .E8(),
    .E9(\net_cnt_lcd_reg[1]_W9_to_E911_7_0 ),
    .E10(),
    .E11(\net_Lut-U196_1_0_W11_to_E1111_7_0 ),
    .E12(),
    .E13(),
    .E14(\net_Lut-U196_1_E14_to_W1411_8_0 ),
    .E15(),
    .E16(\net_Lut-U196_0_1_W16_to_E1611_7_0 ),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(\net_Lut-U205_0_0_S5_to_N511_7_0 ),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(\net_Lut-U205_0_0_S10_to_N1011_7_0 ),
    .N11(),
    .N12(),
    .N13(\net_Lut-U197_0_0_S13_to_N1311_7_0 ),
    .N14(),
    .N15(\net_Lut-U201_0_0_S15_to_N1511_7_0 ),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(\net_cnt_lcd_reg[3]_E8_to_W811_7_0 ),
    .W9(),
    .W10(\net_cnt_lcd_reg[4]_E10_to_W1011_7_0 ),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(net_U113_H6W2_to_H6M211_7_0),
    .H6M3(),
    .H6M4(net_U113_H6W4_to_H6M411_7_0),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(net_U113_V6N2_to_V6M28_7_0),
    .V6N3(),
    .V6N4(),
    .V6N5(net_U113_V6N5_to_V6M58_7_0),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U196_0_1_S0_F_B1_to_F111_7_0 ),
    .S0_F_B2(\net_Lut-U196_1_0_S0_F_B2_to_F211_7_0 ),
    .S0_F_B3(\net_Lut-U197_0_0_S0_F_B3_to_F311_7_0 ),
    .S0_F_B4(\net_Lut-U196_2_1_S0_F_B4_to_F411_7_0 ),
    .S0_G_B1(\net_Lut-U196_3_0_S0_G_B1_to_G111_7_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[4]_S0_G_B2_to_G211_7_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[3]_S0_G_B3_to_G311_7_0 ),
    .S0_G_B4(\net_cnt_lcd_reg[1]_S0_G_B4_to_G411_7_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U196_1_X_to_S0_X11_7_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U196_3_1_Y_to_S0_Y11_7_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U205_0_0_S1_F_B1_to_F111_7_0 ),
    .S1_F_B2(\net_Lut-U204_0_1_S1_F_B2_to_F211_7_0 ),
    .S1_F_B3(\net_cnt_lcd_reg[4]_S1_F_B3_to_F311_7_0 ),
    .S1_F_B4(\net_Lut-U201_0_0_S1_F_B4_to_F411_7_0 ),
    .S1_G_B1(\net_Lut-U205_0_0_S1_G_B1_to_G111_7_0 ),
    .S1_G_B2(\net_Lut-U204_0_1_S1_G_B2_to_G211_7_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[4]_S1_G_B3_to_G311_7_0 ),
    .S1_G_B4(\net_Lut-U201_0_0_S1_G_B4_to_G411_7_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U196_2_1_X_to_S1_X11_7_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U196_3_0_Y_to_S1_Y11_7_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_7_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_7_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_7_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_7_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_7_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_7_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_7_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_7_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_7_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_7_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_7_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_7_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_7_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_7_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_7_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_7_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_7_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_7_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_7_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_7_2_0_inst.sps_v6s2.CONF = "00111101";
  defparam GSB_LFT_7_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_7_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_7_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_7_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_7_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_7_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_7_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_7_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_7_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_7_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_7_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_7_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_7_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_7_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_7_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_7_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(\net_Lut-U126_1_H6W10_to_LEFT_H6E107_2_0 ),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(\net_Lut-U232_0_0_LEFT_H6B7_to_H6M77_3_0 ),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(\net_cnt_lcd_reg[1]_H6W0_to_LEFT_H6M07_2_0 ),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(\net_Lut-U232_0_0_H6W6_to_LEFT_H6M67_2_0 ),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(\net_Lut-U126_1_LEFT_H6D11_to_H6W117_3_0 ),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(\net_cnt_lcd_reg[1]_LEFT_V6S2_to_LEFT_V6M210_2_0 ),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_LFT_10_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_10_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_10_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_10_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_10_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a11.CONF = "110111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_10_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_10_2_0_inst.sps_o1.CONF = "110001101";
  defparam GSB_LFT_10_2_0_inst.sps_o2.CONF = "110101110";
  defparam GSB_LFT_10_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_10_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_10_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_10_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(\net_lcd_db_reg[3]_W15_to_LEFT_E1510_2_0 ),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(\net_lcd_db_reg[4]_W10_to_LEFT_E1010_2_0 ),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(\net_Lut-U157_1_H6W10_to_LEFT_H6E1010_2_0 ),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(\net_cnt_lcd_reg[1]_LEFT_H6A11_to_H6W1110_7_0 ),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(\net_Lut-U157_1_LEFT_H6D11_to_H6W1110_3_0 ),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(\net_cnt_lcd_reg[1]_LEFT_V6S2_to_LEFT_V6M210_2_0 ),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_lcd_db_reg[4]_LEFT_O1_to_OUT10_2_0 ),
    .LEFT_O2(\net_lcd_db_reg[3]_LEFT_O2_to_OUT10_2_0 ),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_10_7_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e12.CONF = "10";
  defparam GSB_CNT_10_7_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_e17.CONF = "10";
  defparam GSB_CNT_10_7_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_e7.CONF = "0";
  defparam GSB_CNT_10_7_0_inst.sps_e8.CONF = "0";
  defparam GSB_CNT_10_7_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_h6e1.CONF = "0010";
  defparam GSB_CNT_10_7_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_7_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_7_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n10.CONF = "10";
  defparam GSB_CNT_10_7_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_n16.CONF = "10";
  defparam GSB_CNT_10_7_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_n20.CONF = "10";
  defparam GSB_CNT_10_7_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_out0.CONF = "000111";
  defparam GSB_CNT_10_7_0_inst.sps_out1.CONF = "001011";
  defparam GSB_CNT_10_7_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_10_7_0_inst.sps_out4.CONF = "011110";
  defparam GSB_CNT_10_7_0_inst.sps_out5.CONF = "011110";
  defparam GSB_CNT_10_7_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s0_f_b1.CONF = "010101111";
  defparam GSB_CNT_10_7_0_inst.sps_s0_f_b2.CONF = "001110111";
  defparam GSB_CNT_10_7_0_inst.sps_s0_f_b3.CONF = "001111011";
  defparam GSB_CNT_10_7_0_inst.sps_s0_f_b4.CONF = "100011111";
  defparam GSB_CNT_10_7_0_inst.sps_s0_g_b1.CONF = "001100";
  defparam GSB_CNT_10_7_0_inst.sps_s0_g_b2.CONF = "011011";
  defparam GSB_CNT_10_7_0_inst.sps_s0_g_b3.CONF = "001011";
  defparam GSB_CNT_10_7_0_inst.sps_s0_g_b4.CONF = "010000";
  defparam GSB_CNT_10_7_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_s13.CONF = "10";
  defparam GSB_CNT_10_7_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s1_f_b1.CONF = "100011111";
  defparam GSB_CNT_10_7_0_inst.sps_s1_f_b2.CONF = "100111101";
  defparam GSB_CNT_10_7_0_inst.sps_s1_f_b3.CONF = "100110111";
  defparam GSB_CNT_10_7_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_7_0_inst.sps_s1_g_b1.CONF = "011010";
  defparam GSB_CNT_10_7_0_inst.sps_s1_g_b2.CONF = "001011";
  defparam GSB_CNT_10_7_0_inst.sps_s1_g_b3.CONF = "001011";
  defparam GSB_CNT_10_7_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_s9.CONF = "0";
  defparam GSB_CNT_10_7_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_7_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_7_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_7_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.sps_w8.CONF = "01";
  defparam GSB_CNT_10_7_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_7_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e0_w0.CONF = "0";
  defparam GSB_CNT_10_7_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n1_e1.CONF = "0";
  defparam GSB_CNT_10_7_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s10_w8.CONF = "0";
  defparam GSB_CNT_10_7_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s15_e13.CONF = "0";
  defparam GSB_CNT_10_7_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s5_e7.CONF = "0";
  defparam GSB_CNT_10_7_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_7_0_inst.switch_s9_w15.CONF = "0";
  GSB_CNT GSB_CNT_10_7_0_inst (
    .E0(\net_cnt_lcd_reg[5]_E0_to_W010_8_0 ),
    .E1(),
    .E2(),
    .E3(\net_Lut-U201_0_0_W3_to_E310_7_0 ),
    .E4(),
    .E5(),
    .E6(\net_cnt_lcd_reg[1]_W6_to_E610_7_0 ),
    .E7(\net_Lut-U205_0_0_E7_to_W710_8_0 ),
    .E8(\net_Lut-U159_0_0_E8_to_W810_8_0 ),
    .E9(),
    .E10(),
    .E11(),
    .E12(\net_Lut-U205_0_0_E12_to_W1210_8_0 ),
    .E13(\net_Lut-U201_0_0_W13_to_E1310_7_0 ),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(\net_Lut-U230_0_0_W20_to_E2010_7_0 ),
    .E21(\net_cnt_lcd_reg[3]_W21_to_E2110_7_0 ),
    .E22(),
    .E23(),
    .N0(),
    .N1(\net_cnt_lcd_reg[4]_S1_to_N110_7_0 ),
    .N2(),
    .N3(\net_cnt_lcd_reg[4]_S3_to_N310_7_0 ),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(\net_Lut-U225_0_N10_to_S109_7_0 ),
    .N11(),
    .N12(\net_Lut-U182_0_1_S12_to_N1210_7_0 ),
    .N13(),
    .N14(),
    .N15(),
    .N16(\net_Lut-U225_0_N16_to_S169_7_0 ),
    .N17(),
    .N18(),
    .N19(),
    .N20(\net_cnt_lcd_reg[1]_N20_to_S209_7_0 ),
    .N21(),
    .N22(),
    .N23(),
    .W0(\net_cnt_lcd_reg[5]_E0_to_W010_7_0 ),
    .W1(\net_cnt_lcd_reg[2]_E1_to_W110_7_0 ),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(\net_cnt_lcd_reg[4]_E10_to_W1010_7_0 ),
    .W11(),
    .W12(\net_Lut-U232_0_0_E12_to_W1210_7_0 ),
    .W13(),
    .W14(),
    .W15(\net_Lut-U225_0_W15_to_E1510_6_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(\net_cnt_lcd_reg[7]_E21_to_W2110_7_0 ),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(\net_Lut-U205_0_0_S5_to_N511_7_0 ),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(\net_Lut-U205_0_0_S10_to_N1011_7_0 ),
    .S11(),
    .S12(),
    .S13(\net_Lut-U197_0_0_S13_to_N1311_7_0 ),
    .S14(),
    .S15(\net_Lut-U201_0_0_S15_to_N1511_7_0 ),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(\net_Lut-U205_0_0_H6E1_to_H6M110_10_0 ),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(\net_Lut-U225_0_H6W1_to_H6M110_7_0 ),
    .H6M2(\net_Lut-U225_0_H6W2_to_H6M210_7_0 ),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(\net_cnt_lcd_reg[1]_LEFT_H6A11_to_H6W1110_7_0 ),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(\net_Lut-U196_6_1_OUT0_to_OUT_W010_8_0 ),
    .OUT1(\net_Lut-U196_7_1_OUT1_to_OUT_W110_8_0 ),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_Lut-U205_0_0_V6S1_to_V6M110_7_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(\net_Lut-U205_0_0_V6S6_to_V6M610_7_0 ),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[7]_S0_F_B1_to_F110_7_0 ),
    .S0_F_B2(\net_Lut-U232_0_0_S0_F_B2_to_F210_7_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[4]_S0_F_B3_to_F310_7_0 ),
    .S0_F_B4(\net_cnt_lcd_reg[2]_S0_F_B4_to_F410_7_0 ),
    .S0_G_B1(\net_Lut-U230_0_0_S0_G_B1_to_G110_7_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[4]_S0_G_B2_to_G210_7_0 ),
    .S0_G_B3(\net_Lut-U201_0_0_S0_G_B3_to_G310_7_0 ),
    .S0_G_B4(\net_Lut-U197_0_0_S0_G_B4_to_G410_7_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U196_6_1_X_to_S0_X10_7_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U196_7_1_Y_to_S0_Y10_7_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[4]_S1_F_B1_to_F110_7_0 ),
    .S1_F_B2(\net_Lut-U201_0_0_S1_F_B2_to_F210_7_0 ),
    .S1_F_B3(\net_Lut-U182_0_1_S1_F_B3_to_F310_7_0 ),
    .S1_F_B4(),
    .S1_G_B1(\net_cnt_lcd_reg[4]_S1_G_B1_to_G110_7_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[3]_S1_G_B2_to_G210_7_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[1]_S1_G_B3_to_G310_7_0 ),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U159_0_0_X_to_S1_X10_7_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U197_0_0_Y_to_S1_Y10_7_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_7_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_e8.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_h6e9.CONF = "001";
  defparam GSB_CNT_9_7_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_7_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_7_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_n15.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_out2.CONF = "001011";
  defparam GSB_CNT_9_7_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_9_7_0_inst.sps_out4.CONF = "011110";
  defparam GSB_CNT_9_7_0_inst.sps_out5.CONF = "000111";
  defparam GSB_CNT_9_7_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s0_f_b1.CONF = "010101111";
  defparam GSB_CNT_9_7_0_inst.sps_s0_f_b2.CONF = "010111101";
  defparam GSB_CNT_9_7_0_inst.sps_s0_f_b3.CONF = "010110111";
  defparam GSB_CNT_9_7_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_7_0_inst.sps_s0_g_b1.CONF = "010010";
  defparam GSB_CNT_9_7_0_inst.sps_s0_g_b2.CONF = "011000";
  defparam GSB_CNT_9_7_0_inst.sps_s0_g_b3.CONF = "100111";
  defparam GSB_CNT_9_7_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_s12.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s1_f_b1.CONF = "100111101";
  defparam GSB_CNT_9_7_0_inst.sps_s1_f_b2.CONF = "100101111";
  defparam GSB_CNT_9_7_0_inst.sps_s1_f_b3.CONF = "110111111";
  defparam GSB_CNT_9_7_0_inst.sps_s1_f_b4.CONF = "010110111";
  defparam GSB_CNT_9_7_0_inst.sps_s1_g_b1.CONF = "100010";
  defparam GSB_CNT_9_7_0_inst.sps_s1_g_b2.CONF = "011000";
  defparam GSB_CNT_9_7_0_inst.sps_s1_g_b3.CONF = "010000";
  defparam GSB_CNT_9_7_0_inst.sps_s1_g_b4.CONF = "001111";
  defparam GSB_CNT_9_7_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_7_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_7_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_7_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w19.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_7_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n12_w17.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n1_w2.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n21_e21.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n5_e5.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s10_e4.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s1_w7.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s3_w5.CONF = "0";
  defparam GSB_CNT_9_7_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_7_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_7_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(\net_Lut-U225_0_E4_to_W49_8_0 ),
    .E5(),
    .E6(),
    .E7(),
    .E8(\net_Lut-U165_2_E8_to_W89_8_0 ),
    .E9(),
    .E10(),
    .E11(),
    .E12(\net_Lut-U201_0_0_W12_to_E129_7_0 ),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(\net_Lut-U190_0_1_E21_to_W219_8_0 ),
    .E22(),
    .E23(),
    .N0(),
    .N1(\net_cnt_lcd_reg[2]_N1_to_S18_7_0 ),
    .N2(\net_Lut-U213_0_0_S2_to_N29_7_0 ),
    .N3(),
    .N4(),
    .N5(\net_Lut-U205_0_0_S5_to_N59_7_0 ),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(\net_Lut-U144_0_0_N12_to_S128_7_0 ),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(\net_Lut-U190_0_1_S21_to_N219_7_0 ),
    .N22(),
    .N23(),
    .W0(),
    .W1(\net_cnt_lcd_reg[5]_E1_to_W19_7_0 ),
    .W2(\net_cnt_lcd_reg[2]_E2_to_W29_7_0 ),
    .W3(),
    .W4(),
    .W5(\net_cnt_lcd_reg[4]_E5_to_W59_7_0 ),
    .W6(),
    .W7(\net_cnt_lcd_reg[4]_E7_to_W79_7_0 ),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(\net_cnt_lcd_reg[3]_E15_to_W159_7_0 ),
    .W16(),
    .W17(\net_Lut-U144_0_0_E17_to_W179_7_0 ),
    .W18(),
    .W19(\net_Lut-U115_0_0_W19_to_E199_6_0 ),
    .W20(\net_cnt_lcd_reg[5]_E20_to_W209_7_0 ),
    .W21(\net_cnt_lcd_reg[1]_E21_to_W219_7_0 ),
    .W22(),
    .W23(),
    .S0(),
    .S1(\net_cnt_lcd_reg[4]_S1_to_N110_7_0 ),
    .S2(),
    .S3(\net_cnt_lcd_reg[4]_S3_to_N310_7_0 ),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(\net_Lut-U225_0_N10_to_S109_7_0 ),
    .S11(),
    .S12(\net_Lut-U182_0_1_S12_to_N1210_7_0 ),
    .S13(),
    .S14(),
    .S15(),
    .S16(\net_Lut-U225_0_N16_to_S169_7_0 ),
    .S17(),
    .S18(),
    .S19(),
    .S20(\net_cnt_lcd_reg[1]_N20_to_S209_7_0 ),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(\net_Lut-U211_0_0_H6E9_to_H6M99_10_0 ),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(\net_Lut-U219_0_1_H6W6_to_H6M69_7_0 ),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(\net_Lut-U166_0_OUT0_to_OUT_W09_7_0 ),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[1]_S0_F_B1_to_F19_7_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[5]_S0_F_B2_to_F29_7_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[3]_S0_F_B3_to_F39_7_0 ),
    .S0_F_B4(),
    .S0_G_B1(\net_cnt_lcd_reg[1]_S0_G_B1_to_G19_7_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[2]_S0_G_B2_to_G29_7_0 ),
    .S0_G_B3(\net_Lut-U213_0_0_S0_G_B3_to_G39_7_0 ),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U182_0_1_X_to_S0_X9_7_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U211_0_0_Y_to_S0_Y9_7_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U225_0_S1_F_B1_to_F19_7_0 ),
    .S1_F_B2(\net_Lut-U205_0_0_S1_F_B2_to_F29_7_0 ),
    .S1_F_B3(\net_Lut-U166_0_S1_F_B3_to_F39_7_0 ),
    .S1_F_B4(\net_Lut-U219_0_1_S1_F_B4_to_F49_7_0 ),
    .S1_G_B1(\net_cnt_lcd_reg[5]_S1_G_B1_to_G19_7_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[1]_S1_G_B2_to_G29_7_0 ),
    .S1_G_B3(\net_cnt_lcd_reg[4]_S1_G_B3_to_G39_7_0 ),
    .S1_G_B4(\net_Lut-U201_0_0_S1_G_B4_to_G49_7_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U165_2_X_to_S1_X9_7_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U115_0_0_Y_to_S1_Y9_7_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_9_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_9_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_9_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_out0.CONF = "011101";
  defparam GSB_CNT_11_9_0_inst.sps_out1.CONF = "011110";
  defparam GSB_CNT_11_9_0_inst.sps_out2.CONF = "001011";
  defparam GSB_CNT_11_9_0_inst.sps_out3.CONF = "011110";
  defparam GSB_CNT_11_9_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_out6.CONF = "000111";
  defparam GSB_CNT_11_9_0_inst.sps_out7.CONF = "011110";
  defparam GSB_CNT_11_9_0_inst.sps_s0.CONF = "0";
  defparam GSB_CNT_11_9_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s0_f_b1.CONF = "100011111";
  defparam GSB_CNT_11_9_0_inst.sps_s0_f_b2.CONF = "001110111";
  defparam GSB_CNT_11_9_0_inst.sps_s0_f_b3.CONF = "100111110";
  defparam GSB_CNT_11_9_0_inst.sps_s0_f_b4.CONF = "010011111";
  defparam GSB_CNT_11_9_0_inst.sps_s0_g_b1.CONF = "011111";
  defparam GSB_CNT_11_9_0_inst.sps_s0_g_b2.CONF = "011000";
  defparam GSB_CNT_11_9_0_inst.sps_s0_g_b3.CONF = "010000";
  defparam GSB_CNT_11_9_0_inst.sps_s0_g_b4.CONF = "110111";
  defparam GSB_CNT_11_9_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s1_f_b1.CONF = "001101111";
  defparam GSB_CNT_11_9_0_inst.sps_s1_f_b2.CONF = "011101111";
  defparam GSB_CNT_11_9_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_9_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_9_0_inst.sps_s1_g_b1.CONF = "001010";
  defparam GSB_CNT_11_9_0_inst.sps_s1_g_b2.CONF = "010000";
  defparam GSB_CNT_11_9_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_9_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_v6n9.CONF = "000";
  defparam GSB_CNT_11_9_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_9_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_9_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_w1.CONF = "0";
  defparam GSB_CNT_11_9_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_w13.CONF = "0";
  defparam GSB_CNT_11_9_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w21.CONF = "10";
  defparam GSB_CNT_11_9_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w7.CONF = "0";
  defparam GSB_CNT_11_9_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_9_0_inst.sps_w9.CONF = "10";
  defparam GSB_CNT_11_9_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e0_w0.CONF = "0";
  defparam GSB_CNT_11_9_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n12_w17.CONF = "0";
  defparam GSB_CNT_11_9_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n21_w22.CONF = "0";
  defparam GSB_CNT_11_9_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n2_e22.CONF = "0";
  defparam GSB_CNT_11_9_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n6_e2.CONF = "0";
  defparam GSB_CNT_11_9_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_n9_w10.CONF = "0";
  defparam GSB_CNT_11_9_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_9_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_9_0_inst (
    .E0(),
    .E1(),
    .E2(\net_cnt_lcd_reg[5]_E2_to_W211_10_0 ),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(\net_cnt_lcd_reg[2]_W7_to_E711_9_0 ),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(\net_cnt_lcd_reg[4]_E22_to_W2211_10_0 ),
    .E23(),
    .N0(),
    .N1(),
    .N2(\net_cnt_lcd_reg[4]_S2_to_N211_9_0 ),
    .N3(),
    .N4(\net_cnt_lcd_reg[5]_S4_to_N411_9_0 ),
    .N5(),
    .N6(\net_cnt_lcd_reg[5]_S6_to_N611_9_0 ),
    .N7(),
    .N8(),
    .N9(\net_cnt_lcd_reg[4]_S9_to_N911_9_0 ),
    .N10(),
    .N11(),
    .N12(\net_Lut-U170_0_S12_to_N1211_9_0 ),
    .N13(),
    .N14(),
    .N15(\net_Lut-U230_0_0_S15_to_N1511_9_0 ),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(\net_cnt_lcd_reg[7]_S20_to_N2011_9_0 ),
    .N21(\net_cnt_lcd_reg[5]_S21_to_N2111_9_0 ),
    .N22(),
    .N23(),
    .W0(\net_cnt_lcd_reg[1]_E0_to_W011_9_0 ),
    .W1(\net_Lut-U204_0_1_W1_to_E111_8_0 ),
    .W2(\net_cnt_lcd_reg[1]_E2_to_W211_9_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(\net_Lut-U215_0_0_W7_to_E711_8_0 ),
    .W8(),
    .W9(\net_Lut-U196_5_1_W9_to_E911_8_0 ),
    .W10(\net_cnt_lcd_reg[4]_W10_to_E1011_8_0 ),
    .W11(),
    .W12(\net_Lut-U232_0_0_E12_to_W1211_9_0 ),
    .W13(\net_Lut-U204_0_1_W13_to_E1311_8_0 ),
    .W14(),
    .W15(),
    .W16(),
    .W17(\net_Lut-U170_0_W17_to_E1711_8_0 ),
    .W18(),
    .W19(),
    .W20(),
    .W21(\net_Lut-U196_4_1_W21_to_E2111_8_0 ),
    .W22(\net_cnt_lcd_reg[5]_W22_to_E2211_8_0 ),
    .W23(),
    .S0(),
    .S1(),
    .S2(\net_cnt_lcd_reg[2]_N2_to_S211_9_0 ),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(\net_Lut-U202_0_0_OUT7_to_OUT_E711_8_0 ),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(\net_Lut-U198_0_0_OUT6_to_OUT_E611_9_0 ),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(\net_Lut-U202_0_0_V6N9_to_V6M98_9_0 ),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(\net_Lut-U204_0_1_V6S8_to_V6M811_9_0 ),
    .V6M9(),
    .V6M10(\net_Lut-U204_0_1_V6S10_to_V6M1011_9_0 ),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[7]_S0_F_B1_to_F111_9_0 ),
    .S0_F_B2(\net_Lut-U232_0_0_S0_F_B2_to_F211_9_0 ),
    .S0_F_B3(\net_Lut-U202_0_0_S0_F_B3_to_F311_9_0 ),
    .S0_F_B4(\net_cnt_lcd_reg[2]_S0_F_B4_to_F411_9_0 ),
    .S0_G_B1(\net_Lut-U230_0_0_S0_G_B1_to_G111_9_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G211_9_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[5]_S0_G_B3_to_G311_9_0 ),
    .S0_G_B4(\net_Lut-U198_0_0_S0_G_B4_to_G411_9_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U196_4_1_X_to_S0_X11_9_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U196_5_1_Y_to_S0_Y11_9_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[1]_S1_F_B1_to_F111_9_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[2]_S1_F_B2_to_F211_9_0 ),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(\net_cnt_lcd_reg[1]_S1_G_B1_to_G111_9_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[5]_S1_G_B2_to_G211_9_0 ),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U215_0_0_X_to_S1_X11_9_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U202_0_0_Y_to_S1_Y11_9_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_h6w10.CONF = "000";
  defparam GSB_CNT_9_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_h6w6.CONF = "000";
  defparam GSB_CNT_9_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n17.CONF = "0";
  defparam GSB_CNT_9_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n23.CONF = "0";
  defparam GSB_CNT_9_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_n4.CONF = "10";
  defparam GSB_CNT_9_8_0_inst.sps_n5.CONF = "0";
  defparam GSB_CNT_9_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_out2.CONF = "001011";
  defparam GSB_CNT_9_8_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_out4.CONF = "011110";
  defparam GSB_CNT_9_8_0_inst.sps_out5.CONF = "001011";
  defparam GSB_CNT_9_8_0_inst.sps_out6.CONF = "011101";
  defparam GSB_CNT_9_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s0_f_b1.CONF = "100111101";
  defparam GSB_CNT_9_8_0_inst.sps_s0_f_b2.CONF = "010101111";
  defparam GSB_CNT_9_8_0_inst.sps_s0_f_b3.CONF = "010101111";
  defparam GSB_CNT_9_8_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_8_0_inst.sps_s0_g_b1.CONF = "010010";
  defparam GSB_CNT_9_8_0_inst.sps_s0_g_b2.CONF = "010111";
  defparam GSB_CNT_9_8_0_inst.sps_s0_g_b3.CONF = "001111";
  defparam GSB_CNT_9_8_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_s12.CONF = "0";
  defparam GSB_CNT_9_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s16.CONF = "10";
  defparam GSB_CNT_9_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s1_f_b1.CONF = "110111111";
  defparam GSB_CNT_9_8_0_inst.sps_s1_f_b2.CONF = "010110111";
  defparam GSB_CNT_9_8_0_inst.sps_s1_f_b3.CONF = "100111101";
  defparam GSB_CNT_9_8_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_8_0_inst.sps_s1_g_b1.CONF = "101111";
  defparam GSB_CNT_9_8_0_inst.sps_s1_g_b2.CONF = "100100";
  defparam GSB_CNT_9_8_0_inst.sps_s1_g_b3.CONF = "100101";
  defparam GSB_CNT_9_8_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s7.CONF = "0";
  defparam GSB_CNT_9_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_v6n5.CONF = "010";
  defparam GSB_CNT_9_8_0_inst.sps_v6n7.CONF = "010";
  defparam GSB_CNT_9_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_8_0_inst.sps_v6s4.CONF = "011";
  defparam GSB_CNT_9_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n11_w12.CONF = "0";
  defparam GSB_CNT_9_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n23_e23.CONF = "0";
  defparam GSB_CNT_9_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n5_e5.CONF = "0";
  defparam GSB_CNT_9_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s19_e17.CONF = "0";
  defparam GSB_CNT_9_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_8_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(\net_cnt_lcd_reg[2]_E5_to_W59_9_0 ),
    .E6(),
    .E7(),
    .E8(),
    .E9(\net_Lut-U224_0_1_W9_to_E99_8_0 ),
    .E10(),
    .E11(\net_Lut-U151_0_W11_to_E119_8_0 ),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(\net_Lut-U230_0_0_W17_to_E179_8_0 ),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(\net_cnt_lcd_reg[3]_E23_to_W239_9_0 ),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(\net_cnt_lcd_reg[2]_N4_to_S48_8_0 ),
    .N5(\net_cnt_lcd_reg[2]_N5_to_S58_8_0 ),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(\net_Lut-U201_0_0_S11_to_N119_8_0 ),
    .N12(\net_cnt_lcd_reg[4]_S12_to_N129_8_0 ),
    .N13(),
    .N14(),
    .N15(),
    .N16(\net_Lut-U170_1_S16_to_N169_8_0 ),
    .N17(\net_cnt_lcd_reg[3]_N17_to_S178_8_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(\net_Lut-U225_0_E4_to_W49_8_0 ),
    .W5(),
    .W6(),
    .W7(),
    .W8(\net_Lut-U165_2_E8_to_W89_8_0 ),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_Lut-U201_0_0_W12_to_E129_7_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(\net_Lut-U190_0_1_E21_to_W219_8_0 ),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(\net_cnt_lcd_reg[1]_N5_to_S59_8_0 ),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(\net_Lut-U164_0_0_S12_to_N1210_8_0 ),
    .S13(),
    .S14(),
    .S15(),
    .S16(\net_cnt_lcd_reg[3]_S16_to_N1610_8_0 ),
    .S17(),
    .S18(),
    .S19(\net_Lut-U230_0_0_S19_to_N1910_8_0 ),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(\net_cnt_lcd_reg[2]_H6E0_to_H6M09_8_0 ),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(\net_cnt_lcd_reg[2]_H6E5_to_H6M59_8_0 ),
    .H6M6(),
    .H6M7(\net_cnt_lcd_reg[3]_H6E7_to_H6M79_8_0 ),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(\net_cnt_lcd_reg[3]_H6E11_to_H6M119_8_0 ),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_Lut-U162_1_H6W6_to_H6M69_5_0 ),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(\net_Lut-U150_0_H6W10_to_LEFT_H6E109_2_0 ),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(\net_Lut-U153_0_OUT6_to_OUT_E69_8_0 ),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(\net_cnt_lcd_reg[2]_V6N5_to_V6M56_8_0 ),
    .V6N6(),
    .V6N7(\net_cnt_lcd_reg[3]_V6N7_to_V6M76_8_0 ),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(\net_cnt_lcd_reg[2]_V6S4_to_V6M412_8_0 ),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[1]_S0_F_B1_to_F19_8_0 ),
    .S0_F_B2(\net_Lut-U170_1_S0_F_B2_to_F29_8_0 ),
    .S0_F_B3(\net_Lut-U224_0_1_S0_F_B3_to_F39_8_0 ),
    .S0_F_B4(),
    .S0_G_B1(\net_Lut-U190_0_1_S0_G_B1_to_G19_8_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[4]_S0_G_B2_to_G29_8_0 ),
    .S0_G_B3(\net_Lut-U201_0_0_S0_G_B3_to_G39_8_0 ),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U162_0_0_X_to_S0_X9_8_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U164_0_0_Y_to_S0_Y9_8_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U153_0_S1_F_B1_to_F19_8_0 ),
    .S1_F_B2(\net_Lut-U225_0_S1_F_B2_to_F29_8_0 ),
    .S1_F_B3(\net_Lut-U151_0_S1_F_B3_to_F39_8_0 ),
    .S1_F_B4(),
    .S1_G_B1(\net_Lut-U162_0_0_S1_G_B1_to_G19_8_0 ),
    .S1_G_B2(\net_Lut-U165_2_S1_G_B2_to_G29_8_0 ),
    .S1_G_B3(\net_Lut-U164_0_0_S1_G_B3_to_G39_8_0 ),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U150_0_X_to_S1_X9_8_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U162_1_Y_to_S1_Y9_8_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_h6w0.CONF = "0011";
  defparam GSB_CNT_11_6_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_6_0_inst.sps_n0.CONF = "10";
  defparam GSB_CNT_11_6_0_inst.sps_n1.CONF = "10";
  defparam GSB_CNT_11_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n13.CONF = "10";
  defparam GSB_CNT_11_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_out0.CONF = "000111";
  defparam GSB_CNT_11_6_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_out4.CONF = "001011";
  defparam GSB_CNT_11_6_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s0_f_b1.CONF = "100111011";
  defparam GSB_CNT_11_6_0_inst.sps_s0_f_b2.CONF = "010110111";
  defparam GSB_CNT_11_6_0_inst.sps_s0_f_b3.CONF = "100110111";
  defparam GSB_CNT_11_6_0_inst.sps_s0_f_b4.CONF = "100011111";
  defparam GSB_CNT_11_6_0_inst.sps_s0_g_b1.CONF = "100101";
  defparam GSB_CNT_11_6_0_inst.sps_s0_g_b2.CONF = "001101";
  defparam GSB_CNT_11_6_0_inst.sps_s0_g_b3.CONF = "010000";
  defparam GSB_CNT_11_6_0_inst.sps_s0_g_b4.CONF = "010111";
  defparam GSB_CNT_11_6_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_6_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n14_e10.CONF = "0";
  defparam GSB_CNT_11_6_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s14_e8.CONF = "0";
  defparam GSB_CNT_11_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s7_n7.CONF = "0";
  defparam GSB_CNT_11_6_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_6_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(\net_cnt_lcd_reg[3]_E8_to_W811_7_0 ),
    .E9(),
    .E10(\net_cnt_lcd_reg[4]_E10_to_W1011_7_0 ),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(\net_Lut-U186_0_N0_to_S010_6_0 ),
    .N1(\net_Lut-U124_0_0_N1_to_S110_6_0 ),
    .N2(\net_cnt_lcd_reg[1]_S2_to_N211_6_0 ),
    .N3(),
    .N4(\net_cnt_lcd_reg[5]_S4_to_N411_6_0 ),
    .N5(),
    .N6(),
    .N7(\net_cnt_lcd_reg[1]_S7_to_N711_6_0 ),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(\net_cnt_lcd_reg[3]_S12_to_N1211_6_0 ),
    .N13(\net_Lut-U123_2_0_N13_to_S1310_6_0 ),
    .N14(\net_cnt_lcd_reg[4]_S14_to_N1411_6_0 ),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(\net_cnt_lcd_reg[2]_E1_to_W111_6_0 ),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(\net_cnt_lcd_reg[3]_N8_to_S811_6_0 ),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(\net_cnt_lcd_reg[3]_N14_to_S1411_6_0 ),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(\net_Lut-U186_0_V6S0_to_V6M011_6_0 ),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[4]_S0_F_B1_to_F111_6_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[3]_S0_F_B2_to_F211_6_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[1]_S0_F_B3_to_F311_6_0 ),
    .S0_F_B4(\net_cnt_lcd_reg[2]_S0_F_B4_to_F411_6_0 ),
    .S0_G_B1(\net_cnt_lcd_reg[4]_S0_G_B1_to_G111_6_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[1]_S0_G_B2_to_G211_6_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[5]_S0_G_B3_to_G311_6_0 ),
    .S0_G_B4(\net_cnt_lcd_reg[3]_S0_G_B4_to_G411_6_0 ),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U124_0_0_X_to_S0_X11_6_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U123_2_0_Y_to_S0_Y11_6_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_11_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_11_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_11_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_11_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_11_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_11_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_11_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e2_w2.CONF = "0";
  defparam GSB_CNT_11_11_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n6_e2.CONF = "0";
  defparam GSB_CNT_11_11_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_11_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_11_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(\net_cnt_lcd_reg[1]_S6_to_N611_11_0 ),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(\net_cnt_lcd_reg[1]_W2_to_E211_10_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_10_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_h6w1.CONF = "0010";
  defparam GSB_CNT_11_10_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_h6w2.CONF = "0010";
  defparam GSB_CNT_11_10_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_h6w4.CONF = "000";
  defparam GSB_CNT_11_10_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_h6w8.CONF = "000";
  defparam GSB_CNT_11_10_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_10_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_10_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n13.CONF = "10";
  defparam GSB_CNT_11_10_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_out0.CONF = "011110";
  defparam GSB_CNT_11_10_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_out2.CONF = "011110";
  defparam GSB_CNT_11_10_0_inst.sps_out3.CONF = "011110";
  defparam GSB_CNT_11_10_0_inst.sps_out4.CONF = "000111";
  defparam GSB_CNT_11_10_0_inst.sps_out5.CONF = "011110";
  defparam GSB_CNT_11_10_0_inst.sps_out6.CONF = "001011";
  defparam GSB_CNT_11_10_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_f_b1.CONF = "101111111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_f_b2.CONF = "011101111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_g_b1.CONF = "011100";
  defparam GSB_CNT_11_10_0_inst.sps_s0_g_b2.CONF = "011111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s1_f_b1.CONF = "011101111";
  defparam GSB_CNT_11_10_0_inst.sps_s1_f_b2.CONF = "100111110";
  defparam GSB_CNT_11_10_0_inst.sps_s1_f_b3.CONF = "010110111";
  defparam GSB_CNT_11_10_0_inst.sps_s1_f_b4.CONF = "001111110";
  defparam GSB_CNT_11_10_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_10_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_10_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_10_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_10_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s0_w2.CONF = "0";
  defparam GSB_CNT_11_10_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s1_n1.CONF = "0";
  defparam GSB_CNT_11_10_0_inst.switch_s1_w7.CONF = "0";
  defparam GSB_CNT_11_10_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_10_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_10_0_inst (
    .E0(),
    .E1(),
    .E2(\net_cnt_lcd_reg[1]_W2_to_E211_10_0 ),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(\net_Lut-U216_0_N13_to_S1310_10_0 ),
    .N14(),
    .N15(),
    .N16(),
    .N17(\net_Lut-U217_1_S17_to_N1711_10_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(\net_cnt_lcd_reg[3]_S21_to_N2111_10_0 ),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(\net_cnt_lcd_reg[5]_E2_to_W211_10_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(\net_cnt_lcd_reg[2]_W7_to_E711_9_0 ),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(\net_cnt_lcd_reg[4]_E22_to_W2211_10_0 ),
    .W23(),
    .S0(),
    .S1(\net_cnt_lcd_reg[2]_N1_to_S111_10_0 ),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(net_U113_H6W1_to_H6E111_4_0),
    .H6W2(net_U113_H6W2_to_H6M211_7_0),
    .H6W3(),
    .H6W4(net_U113_H6W4_to_H6M411_7_0),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(net_U113_H6W8_to_H6E811_4_0),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(\net_Lut-U198_0_0_OUT6_to_OUT_E611_9_0 ),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U216_0_0_S0_F_B1_to_F111_10_0 ),
    .S0_F_B2(\net_Lut-U217_1_S0_F_B2_to_F211_10_0 ),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_cnt_lcd_reg[4]_S0_G_B1_to_G111_10_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[3]_S0_G_B2_to_G211_10_0 ),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U216_0_X_to_S0_X11_10_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U198_0_0_Y_to_S0_Y11_10_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[2]_S1_F_B1_to_F111_10_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[5]_S1_F_B2_to_F211_10_0 ),
    .S1_F_B3(\net_cnt_lcd_reg[3]_S1_F_B3_to_F311_10_0 ),
    .S1_F_B4(\net_cnt_lcd_reg[1]_S1_F_B4_to_F411_10_0 ),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U216_0_0_X_to_S1_X11_10_0 ),
    .S1_XB(),
    .S1_Y(net_U113_Y_to_S1_Y11_10_0),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_10_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_h6w3.CONF = "0001";
  defparam GSB_CNT_8_10_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_10_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_10_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_n12.CONF = "01";
  defparam GSB_CNT_8_10_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_n9.CONF = "10";
  defparam GSB_CNT_8_10_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_8_10_0_inst.sps_out4.CONF = "001011";
  defparam GSB_CNT_8_10_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_out6.CONF = "011110";
  defparam GSB_CNT_8_10_0_inst.sps_out7.CONF = "000111";
  defparam GSB_CNT_8_10_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s0_f_b1.CONF = "011111101";
  defparam GSB_CNT_8_10_0_inst.sps_s0_f_b2.CONF = "011111110";
  defparam GSB_CNT_8_10_0_inst.sps_s0_f_b3.CONF = "010111011";
  defparam GSB_CNT_8_10_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_10_0_inst.sps_s0_g_b1.CONF = "011011";
  defparam GSB_CNT_8_10_0_inst.sps_s0_g_b2.CONF = "011000";
  defparam GSB_CNT_8_10_0_inst.sps_s0_g_b3.CONF = "010101";
  defparam GSB_CNT_8_10_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s19.CONF = "0";
  defparam GSB_CNT_8_10_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s1_f_b1.CONF = "010110111";
  defparam GSB_CNT_8_10_0_inst.sps_s1_f_b2.CONF = "010111101";
  defparam GSB_CNT_8_10_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_10_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_10_0_inst.sps_s1_g_b1.CONF = "001101";
  defparam GSB_CNT_8_10_0_inst.sps_s1_g_b2.CONF = "010100";
  defparam GSB_CNT_8_10_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_10_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_10_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_10_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_10_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e13_w13.CONF = "0";
  defparam GSB_CNT_8_10_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n15_w16.CONF = "0";
  defparam GSB_CNT_8_10_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s5_n5.CONF = "0";
  defparam GSB_CNT_8_10_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_10_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_10_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(\net_cnt_lcd_reg[1]_W9_to_E98_10_0 ),
    .E10(),
    .E11(),
    .E12(),
    .E13(\net_cnt_lcd_reg[1]_W13_to_E138_10_0 ),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(\net_cnt_lcd_reg[3]_W22_to_E228_10_0 ),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(\net_Lut-U229_0_S5_to_N58_10_0 ),
    .N6(),
    .N7(\net_cnt_lcd_reg[1]_S7_to_N78_10_0 ),
    .N8(),
    .N9(\net_Lut-U177_0_0_N9_to_S97_10_0 ),
    .N10(),
    .N11(),
    .N12(\net_Lut-U183_0_0_N12_to_S127_10_0 ),
    .N13(),
    .N14(),
    .N15(\net_Lut-U229_0_S15_to_N158_10_0 ),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(\net_cnt_lcd_reg[5]_E0_to_W08_10_0 ),
    .W1(),
    .W2(\net_cnt_lcd_reg[5]_E2_to_W28_10_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(\net_Lut-U229_0_W16_to_E168_9_0 ),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(\net_Lut-U229_0_S5_to_N59_10_0 ),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(\net_cnt_lcd_reg[3]_N15_to_S158_10_0 ),
    .S16(),
    .S17(),
    .S18(),
    .S19(\net_Lut-U226_0_0_S19_to_N199_10_0 ),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(\net_Lut-U188_0_0_H6W3_to_H6M38_7_0 ),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_cnt_lcd_reg[1]_S0_F_B1_to_F18_10_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[5]_S0_F_B2_to_F28_10_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[3]_S0_F_B3_to_F38_10_0 ),
    .S0_F_B4(),
    .S0_G_B1(\net_cnt_lcd_reg[1]_S0_G_B1_to_G18_10_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[5]_S0_G_B2_to_G28_10_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[3]_S0_G_B3_to_G38_10_0 ),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U188_0_0_X_to_S0_X8_10_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U183_0_0_Y_to_S0_Y8_10_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_cnt_lcd_reg[1]_S1_F_B1_to_F18_10_0 ),
    .S1_F_B2(\net_cnt_lcd_reg[5]_S1_F_B2_to_F28_10_0 ),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(\net_cnt_lcd_reg[3]_S1_G_B1_to_G18_10_0 ),
    .S1_G_B2(\net_cnt_lcd_reg[1]_S1_G_B2_to_G28_10_0 ),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U177_0_0_X_to_S1_X8_10_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U226_0_0_Y_to_S1_Y8_10_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_11_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_11_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_11_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_s8.CONF = "10";
  defparam GSB_CNT_8_11_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_11_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_11_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_11_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_11_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n4_w9.CONF = "0";
  defparam GSB_CNT_8_11_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n8_w13.CONF = "0";
  defparam GSB_CNT_8_11_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s20_w22.CONF = "0";
  defparam GSB_CNT_8_11_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_11_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_11_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(\net_cnt_lcd_reg[1]_S4_to_N48_11_0 ),
    .N5(),
    .N6(),
    .N7(),
    .N8(\net_cnt_lcd_reg[1]_S8_to_N88_11_0 ),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(\net_cnt_lcd_reg[1]_W9_to_E98_10_0 ),
    .W10(),
    .W11(),
    .W12(),
    .W13(\net_cnt_lcd_reg[1]_W13_to_E138_10_0 ),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(\net_cnt_lcd_reg[3]_W22_to_E228_10_0 ),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(\net_Lut-U209_0_0_S8_to_N89_11_0 ),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(\net_cnt_lcd_reg[3]_N20_to_S208_11_0 ),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(\net_Lut-U209_0_0_H6E9_to_H6M98_11_0 ),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_12_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e0.CONF = "10";
  defparam GSB_CNT_12_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_12_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_12_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n13.CONF = "01";
  defparam GSB_CNT_12_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_12_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s2.CONF = "0011";
  defparam GSB_CNT_12_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_12_8_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w2.CONF = "0";
  defparam GSB_CNT_12_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_12_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n1_w2.CONF = "0";
  defparam GSB_CNT_12_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_12_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_12_8_0_inst (
    .E0(\net_cnt_lcd_reg[2]_E0_to_W012_9_0 ),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(\net_cnt_lcd_reg[2]_N1_to_S111_8_0 ),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(\net_cnt_lcd_reg[3]_N13_to_S1311_8_0 ),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(\net_cnt_lcd_reg[3]_H6E2_to_H6M212_8_0 ),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(\net_cnt_lcd_reg[2]_V6S4_to_V6M412_8_0 ),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_12_9_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_12_9_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_12_9_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_12_9_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_12_9_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_12_9_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_12_9_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s2_n2.CONF = "0";
  defparam GSB_CNT_12_9_0_inst.switch_s2_w0.CONF = "0";
  defparam GSB_CNT_12_9_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_12_9_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_12_9_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(\net_cnt_lcd_reg[2]_N2_to_S211_9_0 ),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(\net_cnt_lcd_reg[2]_E0_to_W012_9_0 ),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_11_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_e15.CONF = "10";
  defparam GSB_CNT_9_11_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_11_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_11_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_n20.CONF = "10";
  defparam GSB_CNT_9_11_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s18.CONF = "01";
  defparam GSB_CNT_9_11_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s6.CONF = "01";
  defparam GSB_CNT_9_11_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_11_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_v6n11.CONF = "001";
  defparam GSB_CNT_9_11_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_v6n7.CONF = "001";
  defparam GSB_CNT_9_11_0_inst.sps_v6n9.CONF = "001";
  defparam GSB_CNT_9_11_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_v6s10.CONF = "010";
  defparam GSB_CNT_9_11_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_11_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_11_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_11_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e15_w15.CONF = "0";
  defparam GSB_CNT_9_11_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n20_w1.CONF = "0";
  defparam GSB_CNT_9_11_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n8_w13.CONF = "0";
  defparam GSB_CNT_9_11_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_11_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_11_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(\net_Lut-U209_0_0_S8_to_N89_11_0 ),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(\net_cnt_lcd_reg[3]_N20_to_S208_11_0 ),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(\net_cnt_lcd_reg[3]_W1_to_E19_10_0 ),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(\net_Lut-U209_0_0_W13_to_E139_10_0 ),
    .W14(),
    .W15(\net_cnt_lcd_reg[3]_W15_to_E159_10_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(\net_cnt_lcd_reg[2]_S6_to_N610_11_0 ),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(\net_cnt_lcd_reg[3]_S18_to_N1810_11_0 ),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(\net_cnt_lcd_reg[2]_H6E5_to_H6M59_8_0 ),
    .H6W6(),
    .H6W7(\net_cnt_lcd_reg[3]_H6E7_to_H6M79_8_0 ),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(\net_cnt_lcd_reg[3]_H6E11_to_H6M119_8_0 ),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(\net_cnt_lcd_reg[3]_V6N7_to_V6M76_11_0 ),
    .V6N8(),
    .V6N9(\net_cnt_lcd_reg[3]_V6N9_to_V6M96_11_0 ),
    .V6N10(),
    .V6N11(\net_cnt_lcd_reg[2]_V6N11_to_V6M116_11_0 ),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(\net_cnt_lcd_reg[2]_V6S10_to_V6M1012_11_0 ),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_8_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e22.CONF = "01";
  defparam GSB_CNT_6_8_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_8_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_8_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s18.CONF = "10";
  defparam GSB_CNT_6_8_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s4.CONF = "10";
  defparam GSB_CNT_6_8_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_8_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_8_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_8_0_inst.sps_w0.CONF = "0";
  defparam GSB_CNT_6_8_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w12.CONF = "0";
  defparam GSB_CNT_6_8_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_8_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s14_e8.CONF = "0";
  defparam GSB_CNT_6_8_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_8_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_8_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(\net_Lut-U144_0_0_W8_to_E86_8_0 ),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(\net_cnt_lcd_reg[2]_E22_to_W226_9_0 ),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(\net_cnt_lcd_reg[2]_W0_to_E06_7_0 ),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_cnt_lcd_reg[3]_W12_to_E126_7_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(\net_cnt_lcd_reg[3]_S4_to_N47_8_0 ),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(\net_Lut-U144_0_0_S14_to_N147_8_0 ),
    .S15(),
    .S16(),
    .S17(),
    .S18(\net_cnt_lcd_reg[3]_S18_to_N187_8_0 ),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(\net_cnt_lcd_reg[3]_H6E2_to_H6M26_8_0 ),
    .H6M3(),
    .H6M4(),
    .H6M5(\net_cnt_lcd_reg[3]_H6E5_to_H6M56_8_0 ),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(\net_cnt_lcd_reg[2]_V6N5_to_V6M56_8_0 ),
    .V6M6(),
    .V6M7(\net_cnt_lcd_reg[3]_V6N7_to_V6M76_8_0 ),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_9_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_9_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_9_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_9_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_9_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.sps_w8.CONF = "01";
  defparam GSB_CNT_6_9_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_9_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s20_w22.CONF = "0";
  defparam GSB_CNT_6_9_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_9_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_9_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(\net_Lut-U144_0_0_W8_to_E86_8_0 ),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(\net_cnt_lcd_reg[2]_E22_to_W226_9_0 ),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(\net_cnt_lcd_reg[2]_S20_to_N207_9_0 ),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_Lut-U144_0_0_V6N1_to_V6M16_9_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_7_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_7_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_7_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_7_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_7_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_7_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_7_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s11_w13.CONF = "0";
  defparam GSB_CNT_6_7_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s18_e12.CONF = "0";
  defparam GSB_CNT_6_7_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s6_e0.CONF = "0";
  defparam GSB_CNT_6_7_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s8_w10.CONF = "0";
  defparam GSB_CNT_6_7_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_7_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_7_0_inst (
    .E0(\net_cnt_lcd_reg[2]_W0_to_E06_7_0 ),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(\net_cnt_lcd_reg[3]_W12_to_E126_7_0 ),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(\net_Lut-U144_0_0_E10_to_W106_7_0 ),
    .W11(),
    .W12(),
    .W13(\net_cnt_lcd_reg[3]_E13_to_W136_7_0 ),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(\net_cnt_lcd_reg[2]_S6_to_N67_7_0 ),
    .S7(),
    .S8(\net_Lut-U144_0_0_S8_to_N87_7_0 ),
    .S9(),
    .S10(),
    .S11(\net_cnt_lcd_reg[3]_S11_to_N117_7_0 ),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(\net_cnt_lcd_reg[3]_S18_to_N187_7_0 ),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n1_e1.CONF = "0";
  defparam GSB_CNT_11_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_5_0_inst (
    .E0(),
    .E1(\net_cnt_lcd_reg[2]_E1_to_W111_6_0 ),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(\net_cnt_lcd_reg[2]_S1_to_N111_5_0 ),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_10_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_h6w1.CONF = "0010";
  defparam GSB_CNT_9_10_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_h6w6.CONF = "000";
  defparam GSB_CNT_9_10_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_10_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_10_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n11.CONF = "0";
  defparam GSB_CNT_9_10_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_out2.CONF = "000111";
  defparam GSB_CNT_9_10_0_inst.sps_out3.CONF = "011101";
  defparam GSB_CNT_9_10_0_inst.sps_out4.CONF = "001011";
  defparam GSB_CNT_9_10_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_out6.CONF = "011110";
  defparam GSB_CNT_9_10_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s0_f_b1.CONF = "011111011";
  defparam GSB_CNT_9_10_0_inst.sps_s0_f_b2.CONF = "010111011";
  defparam GSB_CNT_9_10_0_inst.sps_s0_f_b3.CONF = "001111011";
  defparam GSB_CNT_9_10_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_10_0_inst.sps_s0_g_b1.CONF = "100000";
  defparam GSB_CNT_9_10_0_inst.sps_s0_g_b2.CONF = "010101";
  defparam GSB_CNT_9_10_0_inst.sps_s0_g_b3.CONF = "001101";
  defparam GSB_CNT_9_10_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s17.CONF = "10";
  defparam GSB_CNT_9_10_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s1_f_b1.CONF = "100111011";
  defparam GSB_CNT_9_10_0_inst.sps_s1_f_b2.CONF = "100111110";
  defparam GSB_CNT_9_10_0_inst.sps_s1_f_b3.CONF = "100111011";
  defparam GSB_CNT_9_10_0_inst.sps_s1_f_b4.CONF = "011110111";
  defparam GSB_CNT_9_10_0_inst.sps_s1_g_b1.CONF = "011000";
  defparam GSB_CNT_9_10_0_inst.sps_s1_g_b2.CONF = "011111";
  defparam GSB_CNT_9_10_0_inst.sps_s1_g_b3.CONF = "100100";
  defparam GSB_CNT_9_10_0_inst.sps_s1_g_b4.CONF = "100111";
  defparam GSB_CNT_9_10_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_s8.CONF = "01";
  defparam GSB_CNT_9_10_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_10_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_10_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_10_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_10_0_inst.sps_w9.CONF = "10";
  defparam GSB_CNT_9_10_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n15_e15.CONF = "0";
  defparam GSB_CNT_9_10_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s10_w8.CONF = "0";
  defparam GSB_CNT_9_10_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_10_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_10_0_inst (
    .E0(),
    .E1(\net_cnt_lcd_reg[3]_W1_to_E19_10_0 ),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(\net_Lut-U209_0_0_W13_to_E139_10_0 ),
    .E14(),
    .E15(\net_cnt_lcd_reg[3]_W15_to_E159_10_0 ),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(\net_Lut-U229_0_S5_to_N59_10_0 ),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(\net_cnt_lcd_reg[3]_N15_to_S158_10_0 ),
    .N16(),
    .N17(),
    .N18(),
    .N19(\net_Lut-U226_0_0_S19_to_N199_10_0 ),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(\net_cnt_lcd_reg[2]_E5_to_W59_10_0 ),
    .W6(),
    .W7(),
    .W8(\net_Lut-U205_0_0_W8_to_E89_9_0 ),
    .W9(\net_Lut-U224_0_1_W9_to_E99_9_0 ),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(\net_Lut-U224_0_0_N0_to_S09_10_0 ),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(\net_Lut-U224_0_0_N6_to_S69_10_0 ),
    .S7(\net_Lut-U227_0_N7_to_S79_10_0 ),
    .S8(\net_Lut-U223_0_S8_to_N810_10_0 ),
    .S9(\net_Lut-U225_0_N9_to_S99_10_0 ),
    .S10(\net_Lut-U205_0_0_N10_to_S109_10_0 ),
    .S11(),
    .S12(),
    .S13(\net_Lut-U216_0_N13_to_S139_10_0 ),
    .S14(),
    .S15(),
    .S16(),
    .S17(\net_Lut-U208_0_S17_to_N1710_10_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(\net_cnt_lcd_reg[5]_N23_to_S239_10_0 ),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(\net_Lut-U211_0_0_H6E9_to_H6M99_10_0 ),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(\net_Lut-U219_0_1_H6W6_to_H6M69_7_0 ),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U224_0_0_S0_F_B1_to_F19_10_0 ),
    .S0_F_B2(\net_cnt_lcd_reg[5]_S0_F_B2_to_F29_10_0 ),
    .S0_F_B3(\net_cnt_lcd_reg[3]_S0_F_B3_to_F39_10_0 ),
    .S0_F_B4(),
    .S0_G_B1(\net_cnt_lcd_reg[2]_S0_G_B1_to_G19_10_0 ),
    .S0_G_B2(\net_cnt_lcd_reg[5]_S0_G_B2_to_G29_10_0 ),
    .S0_G_B3(\net_cnt_lcd_reg[3]_S0_G_B3_to_G39_10_0 ),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(\net_Lut-U224_0_1_X_to_S0_X9_10_0 ),
    .S0_XB(),
    .S0_Y(\net_Lut-U219_0_1_Y_to_S0_Y9_10_0 ),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U229_0_S1_F_B1_to_F19_10_0 ),
    .S1_F_B2(\net_Lut-U224_0_0_S1_F_B2_to_F29_10_0 ),
    .S1_F_B3(\net_Lut-U227_0_S1_F_B3_to_F39_10_0 ),
    .S1_F_B4(\net_Lut-U226_0_0_S1_F_B4_to_F49_10_0 ),
    .S1_G_B1(\net_Lut-U225_0_S1_G_B1_to_G19_10_0 ),
    .S1_G_B2(\net_Lut-U211_0_0_S1_G_B2_to_G29_10_0 ),
    .S1_G_B3(\net_Lut-U209_0_0_S1_G_B3_to_G39_10_0 ),
    .S1_G_B4(\net_Lut-U216_0_S1_G_B4_to_G49_10_0 ),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(\net_Lut-U223_0_X_to_S1_X9_10_0 ),
    .S1_XB(),
    .S1_Y(\net_Lut-U208_0_Y_to_S1_Y9_10_0 ),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e10.CONF = "01";
  defparam GSB_CNT_6_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e13.CONF = "01";
  defparam GSB_CNT_6_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_h6e0.CONF = "0010";
  defparam GSB_CNT_6_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_h6e2.CONF = "0010";
  defparam GSB_CNT_6_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_h6e5.CONF = "011";
  defparam GSB_CNT_6_5_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_h6w8.CONF = "010";
  defparam GSB_CNT_6_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_5_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(net_rst_nInvLut_E10_to_W106_6_0),
    .E11(),
    .E12(),
    .E13(\net_cnt_lcd_reg[3]_E13_to_W136_6_0 ),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(\net_cnt_lcd_reg[2]_H6E0_to_H6W06_11_0 ),
    .H6E1(),
    .H6E2(\net_cnt_lcd_reg[3]_H6E2_to_H6M26_8_0 ),
    .H6E3(),
    .H6E4(),
    .H6E5(\net_cnt_lcd_reg[3]_H6E5_to_H6M56_8_0 ),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(net_rst_nInvLut_H6W8_to_LEFT_H6M86_2_0),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(\net_cnt_lcd_reg[2]_V6N0_to_V6M06_5_0 ),
    .V6M1(),
    .V6M2(\net_cnt_lcd_reg[3]_V6N2_to_V6M26_5_0 ),
    .V6M3(),
    .V6M4(),
    .V6M5(\net_cnt_lcd_reg[3]_V6N5_to_V6M56_5_0 ),
    .V6M6(),
    .V6M7(net_rst_nInvLut_V6N7_to_V6M76_5_0),
    .V6M8(),
    .V6M9(net_rst_nInvLut_V6N9_to_V6M96_5_0),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_11_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_11_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_11_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_11_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n0.CONF = "0011";
  defparam GSB_CNT_6_11_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_11_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w12.CONF = "0";
  defparam GSB_CNT_6_11_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w18.CONF = "01";
  defparam GSB_CNT_6_11_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w4.CONF = "01";
  defparam GSB_CNT_6_11_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w6.CONF = "01";
  defparam GSB_CNT_6_11_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_11_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_11_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_11_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(\net_cnt_lcd_reg[2]_W4_to_E46_10_0 ),
    .W5(),
    .W6(\net_cnt_lcd_reg[3]_W6_to_E66_10_0 ),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_cnt_lcd_reg[3]_W12_to_E126_10_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(\net_cnt_lcd_reg[2]_W18_to_E186_10_0 ),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(\net_cnt_lcd_reg[2]_H6E0_to_H6W06_11_0 ),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(\net_cnt_lcd_reg[3]_V6N7_to_V6M76_11_0 ),
    .V6M8(),
    .V6M9(\net_cnt_lcd_reg[3]_V6N9_to_V6M96_11_0 ),
    .V6M10(),
    .V6M11(\net_cnt_lcd_reg[2]_V6N11_to_V6M116_11_0 ),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_10_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_10_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_10_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_10_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_10_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_10_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_10_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n22_e18.CONF = "0";
  defparam GSB_CNT_6_10_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s10_e4.CONF = "0";
  defparam GSB_CNT_6_10_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s18_e12.CONF = "0";
  defparam GSB_CNT_6_10_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s22_n22.CONF = "0";
  defparam GSB_CNT_6_10_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s8_e6.CONF = "0";
  defparam GSB_CNT_6_10_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_10_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_10_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(\net_cnt_lcd_reg[2]_W4_to_E46_10_0 ),
    .E5(),
    .E6(\net_cnt_lcd_reg[3]_W6_to_E66_10_0 ),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(\net_cnt_lcd_reg[3]_W12_to_E126_10_0 ),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(\net_cnt_lcd_reg[2]_W18_to_E186_10_0 ),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(\net_cnt_lcd_reg[3]_S8_to_N87_10_0 ),
    .S9(),
    .S10(\net_cnt_lcd_reg[2]_S10_to_N107_10_0 ),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(\net_cnt_lcd_reg[3]_S18_to_N187_10_0 ),
    .S19(),
    .S20(),
    .S21(),
    .S22(\net_cnt_lcd_reg[2]_S22_to_N227_10_0 ),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_12_11_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_12_11_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_12_11_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_12_11_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_12_11_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_12_11_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_w1.CONF = "0";
  defparam GSB_CNT_12_11_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_12_11_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_12_11_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_12_11_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(\net_cnt_lcd_reg[2]_W1_to_E112_10_0 ),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(\net_cnt_lcd_reg[2]_V6S10_to_V6M1012_11_0 ),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_12_10_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_12_10_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_12_10_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_12_10_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_12_10_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_12_10_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_12_10_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n1_e1.CONF = "0";
  defparam GSB_CNT_12_10_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_12_10_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_12_10_0_inst (
    .E0(),
    .E1(\net_cnt_lcd_reg[2]_W1_to_E112_10_0 ),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(\net_cnt_lcd_reg[2]_N1_to_S111_10_0 ),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_12_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e13.CONF = "01";
  defparam GSB_CNT_12_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e19.CONF = "0";
  defparam GSB_CNT_12_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_h6e2.CONF = "0010";
  defparam GSB_CNT_12_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_12_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_12_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_12_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_12_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_12_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_12_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_12_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_12_5_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(\net_cnt_lcd_reg[3]_E13_to_W1312_6_0 ),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(\net_cnt_lcd_reg[3]_E19_to_W1912_6_0 ),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(\net_cnt_lcd_reg[3]_H6E2_to_H6M212_8_0 ),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(\net_cnt_lcd_reg[3]_V6S2_to_V6M212_5_0 ),
    .V6M3(\net_cnt_lcd_reg[3]_V6S3_to_V6M312_5_0 ),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_12_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_12_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_12_6_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_12_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_12_6_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_12_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_12_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n14_w19.CONF = "0";
  defparam GSB_CNT_12_6_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n8_w13.CONF = "0";
  defparam GSB_CNT_12_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_12_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_12_6_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(\net_cnt_lcd_reg[3]_N8_to_S811_6_0 ),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(\net_cnt_lcd_reg[3]_N14_to_S1411_6_0 ),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(\net_cnt_lcd_reg[3]_E13_to_W1312_6_0 ),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(\net_cnt_lcd_reg[3]_E19_to_W1912_6_0 ),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_9_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_9_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_9_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_9_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_9_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_9_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_9_2_0_inst.sps_o1.CONF = "110001110";
  defparam GSB_LFT_9_2_0_inst.sps_o2.CONF = "011111111";
  defparam GSB_LFT_9_2_0_inst.sps_o3.CONF = "110010111";
  defparam GSB_LFT_9_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_9_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_9_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(\net_lcd_db_reg[5]_W16_to_LEFT_E169_2_0 ),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(\net_lcd_db_reg[1]_W11_to_LEFT_E119_2_0 ),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(\net_Lut-U150_0_H6W10_to_LEFT_H6E109_2_0 ),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(\net_cnt_lcd_reg[3]_LEFT_H6B7_to_H6W79_6_0 ),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(\net_cnt_lcd_reg[3]_LEFT_H6B11_to_H6W119_6_0 ),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(\net_cnt_lcd_reg[3]_H6W6_to_LEFT_H6M69_2_0 ),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(\net_cnt_lcd_reg[3]_H6W10_to_LEFT_H6M109_2_0 ),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(\net_Lut-U150_0_LEFT_H6D11_to_H6W119_3_0 ),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(\net_lcd_db_reg[6]_OUT7_to_LEFT_OUT_E79_2_0 ),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_lcd_db_reg[1]_LEFT_O1_to_OUT9_2_0 ),
    .LEFT_O2(\net_lcd_db_reg[6]_LEFT_O2_to_OUT9_2_0 ),
    .LEFT_O3(\net_lcd_db_reg[5]_LEFT_O3_to_OUT9_2_0 ),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_6_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e10.CONF = "01";
  defparam GSB_CNT_6_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_6_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_6_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_6_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e13_w13.CONF = "0";
  defparam GSB_CNT_6_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s8_w10.CONF = "0";
  defparam GSB_CNT_6_6_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_6_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(\net_Lut-U144_0_0_E10_to_W106_7_0 ),
    .E11(),
    .E12(),
    .E13(\net_cnt_lcd_reg[3]_E13_to_W136_7_0 ),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(net_rst_nInvLut_E10_to_W106_6_0),
    .W11(),
    .W12(),
    .W13(\net_cnt_lcd_reg[3]_E13_to_W136_6_0 ),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(net_rst_nInvLut_S8_to_N87_6_0),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(\net_Lut-U144_0_0_V6N7_to_V6M76_6_0 ),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_12_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_12_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_12_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_12_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_v6s1.CONF = "0010";
  defparam GSB_CNT_7_12_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_v6s2.CONF = "0010";
  defparam GSB_CNT_7_12_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_12_0_inst.sps_v6s4.CONF = "010";
  defparam GSB_CNT_7_12_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_12_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_12_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_12_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_12_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_cnt_lcd_reg[4]_H6E1_to_H6W17_12_0 ),
    .H6W2(\net_cnt_lcd_reg[7]_H6E2_to_H6M27_9_0 ),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(\net_cnt_lcd_reg[4]_H6E9_to_H6W97_12_0 ),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(\net_cnt_lcd_reg[4]_V6S1_to_V6M110_12_0 ),
    .V6S2(\net_cnt_lcd_reg[7]_V6S2_to_V6M210_12_0 ),
    .V6S3(),
    .V6S4(\net_cnt_lcd_reg[4]_V6S4_to_V6M410_12_0 ),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_12_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_h6w1.CONF = "0011";
  defparam GSB_CNT_10_12_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_h6w4.CONF = "001";
  defparam GSB_CNT_10_12_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_12_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_12_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_12_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_12_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_12_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_w15.CONF = "10";
  defparam GSB_CNT_10_12_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_w2.CONF = "0";
  defparam GSB_CNT_10_12_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_12_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_12_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_12_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(\net_cnt_lcd_reg[4]_W2_to_E210_11_0 ),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(\net_cnt_lcd_reg[7]_W15_to_E1510_11_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_cnt_lcd_reg[4]_H6W1_to_H6M110_9_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(\net_cnt_lcd_reg[4]_H6W4_to_H6M410_9_0 ),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_cnt_lcd_reg[4]_V6S1_to_V6M110_12_0 ),
    .V6M2(\net_cnt_lcd_reg[7]_V6S2_to_V6M210_12_0 ),
    .V6M3(),
    .V6M4(\net_cnt_lcd_reg[4]_V6S4_to_V6M410_12_0 ),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_4_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_h6e1.CONF = "0010";
  defparam GSB_CNT_4_6_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_6_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_v6s2.CONF = "0100";
  defparam GSB_CNT_4_6_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_6_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_6_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_cnt_lcd_reg[4]_V6N1_to_V6M14_6_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(\net_cnt_lcd_reg[4]_V6S2_to_V6N210_6_0 ),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_7_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n17.CONF = "0";
  defparam GSB_CNT_7_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_n20.CONF = "10";
  defparam GSB_CNT_7_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_out2.CONF = "001110";
  defparam GSB_CNT_7_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_out4.CONF = "001101";
  defparam GSB_CNT_7_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_7_3_0_inst.sps_s0_f_b1.CONF = "010110111";
  defparam GSB_CNT_7_3_0_inst.sps_s0_f_b2.CONF = "100111011";
  defparam GSB_CNT_7_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_3_0_inst.sps_s0_g_b1.CONF = "100100";
  defparam GSB_CNT_7_3_0_inst.sps_s0_g_b2.CONF = "100101";
  defparam GSB_CNT_7_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s0_sr_b.CONF = "011011";
  defparam GSB_CNT_7_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_v6n1.CONF = "0001";
  defparam GSB_CNT_7_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_v6s1.CONF = "0011";
  defparam GSB_CNT_7_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_v6s2.CONF = "0000";
  defparam GSB_CNT_7_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(\net_Lut-U173_1_W12_to_E127_3_0 ),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(net_rst_nInvLut_S8_to_N87_3_0),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(\net_Lut-U232_0_0_N17_to_S176_3_0 ),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(net_U113_N10_to_S107_3_0),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(\net_cnt_lcd_reg[4]_H6W1_to_H6M17_3_0 ),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(\net_Lut-U232_0_0_LEFT_H6B7_to_H6M77_3_0 ),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(\net_Lut-U126_1_LEFT_H6D11_to_H6W117_3_0 ),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBB1_to_GCLK17_3_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(\net_lcd_db_reg[0]_V6N1_to_V6M14_3_0 ),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(\net_cnt_lcd_reg[4]_V6S1_to_V6M110_3_0 ),
    .V6S2(\net_lcd_db_reg[3]_V6S2_to_V6M210_3_0 ),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U173_1_S0_F_B1_to_F17_3_0 ),
    .S0_F_B2(net_U113_S0_F_B2_to_F27_3_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Lut-U126_1_S0_G_B1_to_G17_3_0 ),
    .S0_G_B2(net_U113_S0_G_B2_to_G27_3_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK7_3_0 ),
    .S0_SR_B(net_rst_nInvLut_S0_SR_B_to_SR7_3_0),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_lcd_db_reg[3]_XQ_to_S0_XQ7_3_0 ),
    .S0_YQ(\net_lcd_db_reg[0]_YQ_to_S0_YQ7_3_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e1.CONF = "0010";
  defparam GSB_CNT_10_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n20.CONF = "10";
  defparam GSB_CNT_10_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w15.CONF = "10";
  defparam GSB_CNT_10_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_n9_w10.CONF = "0";
  defparam GSB_CNT_10_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s10_n10.CONF = "0";
  defparam GSB_CNT_10_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(\net_lcd_db_reg[4]_S9_to_N910_3_0 ),
    .N10(net_U113_N10_to_S109_3_0),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(\net_Lut-U157_1_N20_to_S209_3_0 ),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(\net_lcd_db_reg[4]_W10_to_LEFT_E1010_2_0 ),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(\net_lcd_db_reg[3]_W15_to_LEFT_E1510_2_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(net_U113_N10_to_S1010_3_0),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(\net_cnt_lcd_reg[4]_H6E1_to_H6W110_9_0 ),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(\net_Lut-U157_1_LEFT_H6D11_to_H6W1110_3_0 ),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_cnt_lcd_reg[4]_V6S1_to_V6M110_3_0 ),
    .V6M2(\net_lcd_db_reg[3]_V6S2_to_V6M210_3_0 ),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_6_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_6_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_6_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n12.CONF = "01";
  defparam GSB_CNT_6_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out3.CONF = "000111";
  defparam GSB_CNT_6_3_0_inst.sps_out4.CONF = "000111";
  defparam GSB_CNT_6_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_s8.CONF = "10";
  defparam GSB_CNT_6_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_6_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_6_3_0_inst.sps_v6s8.CONF = "001";
  defparam GSB_CNT_6_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_6_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n23_w0.CONF = "0";
  defparam GSB_CNT_6_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s17_w23.CONF = "0";
  defparam GSB_CNT_6_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_6_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_6_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(net_U108_N12_to_S125_3_0),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(net_U113_S23_to_N236_3_0),
    .W0(net_U113_W0_to_LEFT_E06_2_0),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(\net_Lut-U232_0_0_W23_to_LEFT_E236_2_0 ),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(net_rst_nInvLut_S8_to_N87_3_0),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(\net_Lut-U232_0_0_N17_to_S176_3_0 ),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(net_rst_nInvLut_LEFT_H6B9_to_H6M96_3_0),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(net_U108_V6S8_to_V6N812_3_0),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(net_U108_X_to_S0_X6_3_0),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_6_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_6_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_6_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_6_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_6_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_6_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_6_2_0_inst.sps_o1.CONF = "110100111";
  defparam GSB_LFT_6_2_0_inst.sps_o2.CONF = "110001110";
  defparam GSB_LFT_6_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_6_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_6_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_6_2_0_inst (
    .LEFT_E23(\net_Lut-U232_0_0_W23_to_LEFT_E236_2_0 ),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(net_U113_W0_to_LEFT_E06_2_0),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(net_rst_nInvLut_LEFT_H6B9_to_H6M96_3_0),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(net_rst_nInvLut_H6W8_to_LEFT_H6M86_2_0),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(net_U113_LEFT_O1_to_OUT6_2_0),
    .LEFT_O2(\net_Lut-U232_0_0_LEFT_O2_to_OUT6_2_0 ),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_11_4_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_4_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_4_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_n6.CONF = "01";
  defparam GSB_CNT_11_4_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_4_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_v6n2.CONF = "0101";
  defparam GSB_CNT_11_4_0_inst.sps_v6n3.CONF = "0101";
  defparam GSB_CNT_11_4_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_v6n9.CONF = "100";
  defparam GSB_CNT_11_4_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_4_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_4_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w6.CONF = "10";
  defparam GSB_CNT_11_4_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_4_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_4_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_4_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(net_U113_N6_to_S610_4_0),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(net_U113_W6_to_E611_3_0),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(net_U113_H6W1_to_H6E111_4_0),
    .H6E2(net_U113_H6W2_to_H6M211_7_0),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(net_U113_H6W8_to_H6E811_4_0),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(net_U113_V6N2_to_V6M28_4_0),
    .V6N3(net_U113_V6N3_to_V6M38_4_0),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(net_U113_V6N9_to_V6M98_4_0),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_4_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e13.CONF = "01";
  defparam GSB_CNT_8_4_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e19.CONF = "0";
  defparam GSB_CNT_8_4_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_h6e2.CONF = "0010";
  defparam GSB_CNT_8_4_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_4_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_4_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s16.CONF = "01";
  defparam GSB_CNT_8_4_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_4_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_4_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_4_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_w15.CONF = "10";
  defparam GSB_CNT_8_4_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w6.CONF = "01";
  defparam GSB_CNT_8_4_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_4_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s8_w10.CONF = "0";
  defparam GSB_CNT_8_4_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_4_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_4_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(net_U113_E13_to_W138_5_0),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(net_U113_E19_to_W198_5_0),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(net_U113_W6_to_E68_3_0),
    .W7(),
    .W8(),
    .W9(),
    .W10(\net_lcd_db_reg[2]_W10_to_E108_3_0 ),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(net_U113_W15_to_E158_3_0),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(\net_lcd_db_reg[2]_N8_to_S88_4_0 ),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(net_U113_S16_to_N169_4_0),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(net_U113_V6N2_to_V6M28_4_0),
    .V6M3(net_U113_V6N3_to_V6M38_4_0),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(net_U113_V6N9_to_V6M98_4_0),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_8_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_8_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_8_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_8_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_8_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_8_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e10_w10.CONF = "0";
  defparam GSB_CNT_8_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n10_e6.CONF = "0";
  defparam GSB_CNT_8_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s13_e15.CONF = "0";
  defparam GSB_CNT_8_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_8_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_8_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(net_U113_W6_to_E68_3_0),
    .E7(),
    .E8(),
    .E9(),
    .E10(\net_lcd_db_reg[2]_W10_to_E108_3_0 ),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(net_U113_W15_to_E158_3_0),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(net_U113_N10_to_S107_3_0),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(\net_lcd_db_reg[2]_W10_to_LEFT_E108_2_0 ),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(net_U113_S13_to_N139_3_0),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_11_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_11_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_11_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s10.CONF = "01";
  defparam GSB_CNT_11_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_11_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_11_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_11_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n10_e6.CONF = "0";
  defparam GSB_CNT_11_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_11_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_11_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(net_U113_W6_to_E611_3_0),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(net_U113_N10_to_S1010_3_0),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(\net_Buf-pad-rst_n_S10_to_N1012_3_0 ),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(\net_Buf-pad-rst_n_V6S1_to_V6N111_3_0 ),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n20.CONF = "10";
  defparam GSB_CNT_9_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out3.CONF = "100111";
  defparam GSB_CNT_9_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out5.CONF = "001110";
  defparam GSB_CNT_9_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_out7.CONF = "001101";
  defparam GSB_CNT_9_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b1.CONF = "100011111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b2.CONF = "100111011";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b1.CONF = "011100";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b2.CONF = "100101";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s0_sr_b.CONF = "010111";
  defparam GSB_CNT_9_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s11.CONF = "0";
  defparam GSB_CNT_9_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_clk_b.CONF = "101011";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b1.CONF = "011111011";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b2.CONF = "011111101";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_s1_sr_b.CONF = "010111";
  defparam GSB_CNT_9_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w11.CONF = "10";
  defparam GSB_CNT_9_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w16.CONF = "10";
  defparam GSB_CNT_9_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s20_w22.CONF = "0";
  defparam GSB_CNT_9_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s9_e11.CONF = "0";
  defparam GSB_CNT_9_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(net_rst_nInvLut_W10_to_E109_3_0),
    .E11(\net_lcd_db_reg[4]_W11_to_E119_3_0 ),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(net_U113_S13_to_N139_3_0),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(\net_lcd_db_reg[1]_W11_to_LEFT_E119_2_0 ),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(\net_lcd_db_reg[5]_W16_to_LEFT_E169_2_0 ),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(\net_lcd_db_reg[4]_S9_to_N910_3_0 ),
    .S10(net_U113_N10_to_S109_3_0),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(\net_Lut-U157_1_N20_to_S209_3_0 ),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(\net_Lut-U115_1_H6W8_to_H6M89_3_0 ),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(\net_Lut-U150_0_LEFT_H6D11_to_H6W119_3_0 ),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBD1_to_GCLK19_3_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(\net_lcd_db_reg[6]_OUT7_to_LEFT_OUT_E79_2_0 ),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U150_0_S0_F_B1_to_F19_3_0 ),
    .S0_F_B2(net_U113_S0_F_B2_to_F29_3_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Lut-U157_1_S0_G_B1_to_G19_3_0 ),
    .S0_G_B2(net_U113_S0_G_B2_to_G29_3_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK9_3_0 ),
    .S0_SR_B(net_rst_nInvLut_S0_SR_B_to_SR9_3_0),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_lcd_db_reg[6]_XQ_to_S0_XQ9_3_0 ),
    .S0_YQ(\net_lcd_db_reg[5]_YQ_to_S0_YQ9_3_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(\net_Lut-U115_1_S1_F_B1_to_F19_3_0 ),
    .S1_F_B2(net_U113_S1_F_B2_to_F29_3_0),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(\net_IBuf-clkpad-clk_S1_CLK_B_to_CLK9_3_0 ),
    .S1_SR_B(net_rst_nInvLut_S1_SR_B_to_SR9_3_0),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(\net_lcd_db_reg[1]_XQ_to_S1_XQ9_3_0 ),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_9_4_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_9_4_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_9_4_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_n8.CONF = "01";
  defparam GSB_CNT_9_4_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_out2.CONF = "001101";
  defparam GSB_CNT_9_4_0_inst.sps_out3.CONF = "001110";
  defparam GSB_CNT_9_4_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s0_clk_b.CONF = "111011";
  defparam GSB_CNT_9_4_0_inst.sps_s0_f_b1.CONF = "001011111";
  defparam GSB_CNT_9_4_0_inst.sps_s0_f_b2.CONF = "010101111";
  defparam GSB_CNT_9_4_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_4_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_4_0_inst.sps_s0_g_b1.CONF = "010111";
  defparam GSB_CNT_9_4_0_inst.sps_s0_g_b2.CONF = "010010";
  defparam GSB_CNT_9_4_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s0_sr_b.CONF = "010111";
  defparam GSB_CNT_9_4_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_9_4_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_9_4_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_9_4_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w11.CONF = "10";
  defparam GSB_CNT_9_4_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_9_4_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e10_w10.CONF = "0";
  defparam GSB_CNT_9_4_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_9_4_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_9_4_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(net_rst_nInvLut_W10_to_E109_4_0),
    .E11(),
    .E12(\net_Lut-U162_1_W12_to_E129_4_0 ),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(\net_Lut-U195_1_W20_to_E209_4_0 ),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(\net_lcd_db_reg[2]_N8_to_S88_4_0 ),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(net_U113_S16_to_N169_4_0),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(net_rst_nInvLut_W10_to_E109_3_0),
    .W11(\net_lcd_db_reg[4]_W11_to_E119_3_0 ),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBD1_to_GCLK19_3_0 ),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(\net_Lut-U195_1_S0_F_B1_to_F19_4_0 ),
    .S0_F_B2(net_U113_S0_F_B2_to_F29_4_0),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(\net_Lut-U162_1_S0_G_B1_to_G19_4_0 ),
    .S0_G_B2(net_U113_S0_G_B2_to_G29_4_0),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(\net_IBuf-clkpad-clk_S0_CLK_B_to_CLK9_4_0 ),
    .S0_SR_B(net_rst_nInvLut_S0_SR_B_to_SR9_4_0),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(\net_lcd_db_reg[2]_XQ_to_S0_XQ9_4_0 ),
    .S0_YQ(\net_lcd_db_reg[4]_YQ_to_S0_YQ9_4_0 ),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_10_4_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_10_4_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_10_4_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_10_4_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_10_4_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_10_4_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_10_4_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s6_e0.CONF = "0";
  defparam GSB_CNT_10_4_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_10_4_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_10_4_0_inst (
    .E0(net_U113_E0_to_W010_5_0),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(net_U113_N6_to_S610_4_0),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_4_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_4_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_4_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_4_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_4_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_4_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w21.CONF = "01";
  defparam GSB_CNT_5_4_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_4_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_4_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_4_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(net_U113_W21_to_E215_3_0),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(net_U113_V6N3_to_V6M38_4_0),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s1.CONF = "0011";
  defparam GSB_CNT_5_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s12_w14.CONF = "0";
  defparam GSB_CNT_5_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s23_e21.CONF = "0";
  defparam GSB_CNT_5_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(net_U113_W21_to_E215_3_0),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(net_U108_W14_to_LEFT_E145_2_0),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(net_U108_N12_to_S125_3_0),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(net_U113_S23_to_N236_3_0),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(\net_Buf-pad-rst_n_H6W1_to_H6M15_3_0 ),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(\net_Buf-pad-rst_n_V6S1_to_V6N111_3_0 ),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_RHT_5_54_0_inst.sps_h6w0.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w10.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w4.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w6.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6w8.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_llh0.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh6.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_RHT_5_54_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_RHT_5_54_0_inst.sps_out6.CONF = "1111";
  defparam GSB_RHT_5_54_0_inst.sps_out7.CONF = "1111";
  defparam GSB_RHT_5_54_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_w0.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w1.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w10.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w11.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w12.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w13.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w14.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w15.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w16.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w17.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w18.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w19.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w2.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w20.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w21.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w22.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w23.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w3.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w4.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w5.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w6.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.sps_w7.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w8.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_w9.CONF = "111";
  defparam GSB_RHT_5_54_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_RHT_5_54_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_RHT_5_54_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_llh1.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh10.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh11.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh2.CONF = "01";
  defparam GSB_RHT_5_54_0_inst.sps_llh3.CONF = "01";
  defparam GSB_RHT_5_54_0_inst.sps_llh4.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh5.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh7.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh8.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_llh9.CONF = "11";
  defparam GSB_RHT_5_54_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_RHT_5_54_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_RHT_5_54_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_RHT_5_54_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d10.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d4.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d6.CONF = "111111";
  defparam GSB_RHT_5_54_0_inst.sps_h6d8.CONF = "111111";
  GSB_RHT GSB_RHT_5_54_0_inst (
    .RIGHT_W23(),
    .RIGHT_W22(),
    .RIGHT_W21(),
    .RIGHT_W20(),
    .RIGHT_W19(),
    .RIGHT_W18(),
    .RIGHT_W17(),
    .RIGHT_W16(),
    .RIGHT_W15(),
    .RIGHT_W14(),
    .RIGHT_W13(),
    .RIGHT_W12(),
    .RIGHT_W11(),
    .RIGHT_W10(),
    .RIGHT_W9(),
    .RIGHT_W8(),
    .RIGHT_W7(),
    .RIGHT_W6(),
    .RIGHT_W5(),
    .RIGHT_W4(),
    .RIGHT_W3(),
    .RIGHT_W2(),
    .RIGHT_W1(),
    .RIGHT_W0(),
    .RIGHT_H6A0(),
    .RIGHT_H6A1(),
    .RIGHT_H6A2(),
    .RIGHT_H6A3(),
    .RIGHT_H6A4(),
    .RIGHT_H6A5(),
    .RIGHT_H6A6(),
    .RIGHT_H6A7(),
    .RIGHT_H6A8(),
    .RIGHT_H6A9(),
    .RIGHT_H6A10(),
    .RIGHT_H6A11(),
    .RIGHT_H6B0(),
    .RIGHT_H6B1(),
    .RIGHT_H6B2(),
    .RIGHT_H6B3(),
    .RIGHT_H6B4(),
    .RIGHT_H6B5(),
    .RIGHT_H6B6(),
    .RIGHT_H6B7(),
    .RIGHT_H6B8(),
    .RIGHT_H6B9(),
    .RIGHT_H6B10(),
    .RIGHT_H6B11(),
    .RIGHT_H6M0(),
    .RIGHT_H6M1(),
    .RIGHT_H6M2(),
    .RIGHT_H6M3(),
    .RIGHT_H6M4(),
    .RIGHT_H6M5(),
    .RIGHT_H6M6(),
    .RIGHT_H6M7(),
    .RIGHT_H6M8(),
    .RIGHT_H6M9(),
    .RIGHT_H6M10(),
    .RIGHT_H6M11(),
    .RIGHT_H6C0(),
    .RIGHT_H6C1(),
    .RIGHT_H6C2(),
    .RIGHT_H6C3(),
    .RIGHT_H6C4(),
    .RIGHT_H6C5(),
    .RIGHT_H6C6(),
    .RIGHT_H6C7(),
    .RIGHT_H6C8(),
    .RIGHT_H6C9(),
    .RIGHT_H6C10(),
    .RIGHT_H6C11(),
    .RIGHT_H6D0(),
    .RIGHT_H6D1(),
    .RIGHT_H6D2(),
    .RIGHT_H6D3(),
    .RIGHT_H6D4(),
    .RIGHT_H6D5(),
    .RIGHT_H6D6(),
    .RIGHT_H6D7(),
    .RIGHT_H6D8(),
    .RIGHT_H6D9(),
    .RIGHT_H6D10(),
    .RIGHT_H6D11(),
    .RIGHT_H6W0(),
    .RIGHT_H6W1(),
    .RIGHT_H6W2(),
    .RIGHT_H6W3(),
    .RIGHT_H6W4(),
    .RIGHT_H6W5(),
    .RIGHT_H6W6(),
    .RIGHT_H6W7(),
    .RIGHT_H6W8(),
    .RIGHT_H6W9(),
    .RIGHT_H6W10(),
    .RIGHT_H6W11(),
    .RIGHT_LLH0(),
    .RIGHT_LLH1(),
    .RIGHT_LLH2(\net_Buf-pad-rst_n_RIGHT_LLH2_to_LLH05_5_0 ),
    .RIGHT_LLH3(\net_Buf-pad-rst_n_RIGHT_LLH3_to_LLH05_6_0 ),
    .RIGHT_LLH4(),
    .RIGHT_LLH5(),
    .RIGHT_LLH6(),
    .RIGHT_LLH7(),
    .RIGHT_LLH8(),
    .RIGHT_LLH9(),
    .RIGHT_LLH10(),
    .RIGHT_LLH11(),
    .RIGHT_GCLK0(),
    .RIGHT_GCLK1(),
    .RIGHT_GCLK2(),
    .RIGHT_GCLK3(),
    .RIGHT_OUT_W0(),
    .RIGHT_OUT_W1(),
    .RIGHT_OUT6(),
    .RIGHT_OUT7(),
    .RIGHT_TBUFO2(),
    .RIGHT_TBUFO3(),
    .RIGHT_TBUFO0(),
    .RIGHT_TBUFO1(),
    .RIGHT_V6N0(),
    .RIGHT_V6N1(),
    .RIGHT_V6N2(),
    .RIGHT_V6N3(),
    .RIGHT_V6A0(),
    .RIGHT_V6A1(),
    .RIGHT_V6A2(),
    .RIGHT_V6A3(),
    .RIGHT_V6B0(),
    .RIGHT_V6B1(),
    .RIGHT_V6B2(),
    .RIGHT_V6B3(),
    .RIGHT_V6M0(),
    .RIGHT_V6M1(),
    .RIGHT_V6M2(),
    .RIGHT_V6M3(),
    .RIGHT_V6C0(),
    .RIGHT_V6C1(),
    .RIGHT_V6C2(),
    .RIGHT_V6C3(),
    .RIGHT_V6D0(),
    .RIGHT_V6D1(),
    .RIGHT_V6D2(),
    .RIGHT_V6D3(),
    .RIGHT_V6S0(),
    .RIGHT_V6S1(),
    .RIGHT_V6S2(),
    .RIGHT_V6S3(),
    .RIGHT_LLV0(),
    .RIGHT_LLV6(),
    .RIGHT_PCI_CE(),
    .RIGHT_I1(),
    .RIGHT_I2(),
    .RIGHT_I3(\net_Buf-pad-rst_n_IN_to_RIGHT_I35_54_0 ),
    .RIGHT_IQ1(),
    .RIGHT_IQ2(),
    .RIGHT_IQ3(),
    .RIGHT_ICE1(),
    .RIGHT_ICE2(),
    .RIGHT_ICE3(),
    .RIGHT_O1(),
    .RIGHT_O2(),
    .RIGHT_O3(),
    .RIGHT_OCE1(),
    .RIGHT_OCE2(),
    .RIGHT_OCE3(),
    .RIGHT_T1(),
    .RIGHT_T2(),
    .RIGHT_T3(),
    .RIGHT_TCE1(),
    .RIGHT_TCE2(),
    .RIGHT_TCE3(),
    .RIGHT_CLK1(),
    .RIGHT_CLK2(),
    .RIGHT_CLK3(),
    .RIGHT_SR_B1(),
    .RIGHT_SR_B2(),
    .RIGHT_SR_B3(),
    .RIGHT_TO0(),
    .RIGHT_TO1(),
    .RIGHT_TI0_B(),
    .RIGHT_TI1_B(),
    .RIGHT_TS0_B(),
    .RIGHT_TS1_B()
  );

  defparam GSB_CNT_5_5_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w1.CONF = "0001";
  defparam GSB_CNT_5_5_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_5_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_5_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_5_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s1.CONF = "0010";
  defparam GSB_CNT_5_5_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_5_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_5_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_5_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_5_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_Buf-pad-rst_n_RIGHT_LLH2_to_LLH05_5_0 ),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(\net_Buf-pad-rst_n_V6S1_to_V6M18_5_0 ),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_5_6_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w1.CONF = "0001";
  defparam GSB_CNT_5_6_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_5_6_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_5_6_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_5_6_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_5_6_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_5_6_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_5_6_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_5_6_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(\net_Buf-pad-rst_n_H6W1_to_H6M15_3_0 ),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(\net_Buf-pad-rst_n_RIGHT_LLH3_to_LLH05_6_0 ),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_12_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_12_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_12_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s5.CONF = "01";
  defparam GSB_CNT_12_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_12_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_12_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_12_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_12_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s10_n10.CONF = "0";
  defparam GSB_CNT_12_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_12_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_12_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(\net_Buf-pad-rst_n_S10_to_N1012_3_0 ),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(net_U108_S5_to_N513_3_0),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(\net_Buf-pad-rst_n_S10_to_N1013_3_0 ),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(net_U108_V6S8_to_V6N812_3_0),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CNT_13_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_13_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_13_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_13_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_13_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_13_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n10_w15.CONF = "0";
  defparam GSB_CNT_13_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s5_n5.CONF = "0";
  defparam GSB_CNT_13_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_13_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_13_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(net_U108_S5_to_N513_3_0),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(\net_Buf-pad-rst_n_S10_to_N1013_3_0 ),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(\net_Buf-pad-rst_n_W15_to_LEFT_E1513_2_0 ),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(net_U108_S5_to_N514_3_0),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_13_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_13_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_13_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_13_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_13_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_13_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_13_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_13_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_13_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_13_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_13_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_13_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_13_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_13_2_0_inst.sps_o3.CONF = "110101110";
  defparam GSB_LFT_13_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_13_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_13_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(\net_Buf-pad-rst_n_W15_to_LEFT_E1513_2_0 ),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(),
    .LEFT_O3(\net_Buf-pad-rst_n_LEFT_O3_to_OUT13_2_0 ),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_7_4_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_7_4_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_7_4_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s14.CONF = "10";
  defparam GSB_CNT_7_4_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_7_4_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_7_4_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_7_4_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_7_4_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s14_w12.CONF = "0";
  defparam GSB_CNT_7_4_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_7_4_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_7_4_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(\net_Lut-U173_1_W12_to_E127_3_0 ),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(\net_Lut-U173_1_H6W6_to_H6M67_4_0 ),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_CLKB_35_28_0_inst.sps_h6e0.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e1.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e2.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6e3.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6d0.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6d1.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6d2.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_h6d3.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh1.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh10.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh4.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_llh7.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.spbu_gclk0.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_gclk1.CONF = "0";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e0.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e1.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e2.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_e3.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w0.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w1.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w2.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.spbu_hgclk_w3.CONF = "1";
  defparam GSB_CLKB_35_28_0_inst.sps_ce0.CONF = "1111";
  defparam GSB_CLKB_35_28_0_inst.sps_ce1.CONF = "1111";
  defparam GSB_CLKB_35_28_0_inst.sps_clkfbl.CONF = "010";
  defparam GSB_CLKB_35_28_0_inst.sps_clkfbr.CONF = "010";
  defparam GSB_CLKB_35_28_0_inst.sps_clkinl.CONF = "011";
  defparam GSB_CLKB_35_28_0_inst.sps_clkinr.CONF = "011";
  defparam GSB_CLKB_35_28_0_inst.sps_gclkbuf0_in.CONF = "111111";
  defparam GSB_CLKB_35_28_0_inst.sps_gclkbuf1_in.CONF = "011111";
  GSB_CLKB GSB_CLKB_35_28_0_inst (
    .CLKB_H6E0(),
    .CLKB_H6E1(),
    .CLKB_H6E2(),
    .CLKB_H6E3(),
    .CLKB_H6A0(),
    .CLKB_H6A1(),
    .CLKB_H6A2(),
    .CLKB_H6A3(),
    .CLKB_H6B0(),
    .CLKB_H6B1(),
    .CLKB_H6B2(),
    .CLKB_H6B3(),
    .CLKB_H6M0(),
    .CLKB_H6M1(),
    .CLKB_H6M2(),
    .CLKB_H6M3(),
    .CLKB_H6C0(),
    .CLKB_H6C1(),
    .CLKB_H6C2(),
    .CLKB_H6C3(),
    .CLKB_H6D0(),
    .CLKB_H6D1(),
    .CLKB_H6D2(),
    .CLKB_H6D3(),
    .CLKB_LLH1(),
    .CLKB_LLH4(),
    .CLKB_LLH7(),
    .CLKB_LLH10(),
    .CLKB_GCLK0(),
    .CLKB_GCLK1(\net_IBuf-clkpad-clk_CLKB_GCLK1_to_CLKC_GCLK118_28_0 ),
    .CLKB_VGCLK0(),
    .CLKB_VGCLK1(),
    .CLKB_VGCLK2(),
    .CLKB_VGCLK3(),
    .CLKB_HGCLK_E0(),
    .CLKB_HGCLK_E1(),
    .CLKB_HGCLK_E2(),
    .CLKB_HGCLK_E3(),
    .CLKB_HGCLK_W0(),
    .CLKB_HGCLK_W1(),
    .CLKB_HGCLK_W2(),
    .CLKB_HGCLK_W3(),
    .CLKB_CLKINL_1(),
    .CLKB_CLKFBL_1(),
    .CLKB_CLKDVL_1(),
    .CLKB_CLK0L_1(),
    .CLKB_CLK90L_1(),
    .CLKB_CLK180L_1(),
    .CLKB_CLK270L_1(),
    .CLKB_CLK2XL_1(),
    .CLKB_CLK2X90L_1(),
    .CLKB_LOCKEDL_1(),
    .CLKB_CLKINR_1(),
    .CLKB_CLKFBR_1(),
    .CLKB_CLKDVR_1(),
    .CLKB_CLK0R_1(),
    .CLKB_CLK90R_1(),
    .CLKB_CLK180R_1(),
    .CLKB_CLK270R_1(),
    .CLKB_CLK2XR_1(),
    .CLKB_CLK2X90R_1(),
    .CLKB_LOCKEDR_1(),
    .CLKB_CLKPAD0(),
    .CLKB_CLKPAD1(\net_Buf-pad-clk_GCLKOUT_to_CLKB_CLKPAD135_28_0 ),
    .CLKB_GCLKBUF0_IN(),
    .CLKB_GCLK0_PW(),
    .CLKB_CE0(),
    .CLKB_GCLKBUF1_IN(\net_Buf-pad-clk_CLKB_GCLKBUF1_IN_to_IN35_28_0 ),
    .CLKB_GCLK1_PW(\net_IBuf-clkpad-clk_OUT_to_CLKB_GCLK1_PW35_28_0 ),
    .CLKB_CE1(),
    .BOT_CLKINL(),
    .BOT_CLKFBL(),
    .BOT_CLKINR(),
    .BOT_CLKFBR(),
    .DLL1_RST_I(),
    .DLL1_RST_O(),
    .DLL0_RST_I(),
    .DLL0_RST_O()
  );

  defparam GSB_CNT_14_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_14_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_14_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_14_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_14_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.sps_w8.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_14_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n5_w6.CONF = "0";
  defparam GSB_CNT_14_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_14_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_14_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(net_U108_S5_to_N514_3_0),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(net_U108_W6_to_LEFT_E614_2_0),
    .W7(),
    .W8(),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_14_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_14_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_14_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_14_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_14_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_14_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_14_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_14_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_14_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_14_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_14_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_14_2_0_inst.sps_o1.CONF = "110011101";
  defparam GSB_LFT_14_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_14_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_14_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_14_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_14_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(net_U108_W6_to_LEFT_E614_2_0),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(net_U108_LEFT_O1_to_OUT14_2_0),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_LFT_5_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_5_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_5_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_5_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_5_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_5_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_5_2_0_inst.sps_o1.CONF = "111111111";
  defparam GSB_LFT_5_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_5_2_0_inst.sps_o3.CONF = "110101101";
  defparam GSB_LFT_5_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_5_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_5_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(net_U108_W14_to_LEFT_E145_2_0),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(),
    .LEFT_O2(),
    .LEFT_O3(net_U108_LEFT_O3_to_OUT5_2_0),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_LFT_8_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_8_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_8_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_8_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_8_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_8_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_8_2_0_inst.sps_o1.CONF = "110001101";
  defparam GSB_LFT_8_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_8_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_8_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_8_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_8_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(\net_lcd_db_reg[2]_W10_to_LEFT_E108_2_0 ),
    .LEFT_E9(),
    .LEFT_E8(),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_lcd_db_reg[2]_LEFT_O1_to_OUT8_2_0 ),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  defparam GSB_CNT_4_3_0_inst.spbu_tbuf0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.spbu_tbuf3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e0.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e1.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e11.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e12.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e13.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e15.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e17.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e21.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e23.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e3.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e5.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_e7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_e9.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_h6e0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e11.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e5.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e7.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6e9.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w10.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w4.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w6.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_h6w8.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_llh0.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_llh6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_llv0.CONF = "11111";
  defparam GSB_CNT_4_3_0_inst.sps_llv6.CONF = "11111";
  defparam GSB_CNT_4_3_0_inst.sps_n0.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n1.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n12.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n13.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n16.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n19.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n20.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n21.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n4.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_n6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n7.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n8.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_n9.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_out0.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out2.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out3.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out4.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out5.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out6.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_out7.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s0_bx_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_by_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_ce_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_clk_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b2.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b3.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_g_b4.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s0_sr_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s13.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s14.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s15.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s16.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s17.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s1_bx_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_by_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_ce_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_clk_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b1.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b2.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b3.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_f_b4.CONF = "111111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b2.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b3.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_g_b4.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s1_sr_b.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_s2.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s20.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s3.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s4.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s5.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_s8.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_s9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_ts_b0.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_ts_b1.CONF = "111111";
  defparam GSB_CNT_4_3_0_inst.sps_t_in0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_t_in1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n11.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n5.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n7.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6n9.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s0.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s1.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s10.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s2.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s3.CONF = "1111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s4.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s6.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_v6s8.CONF = "111";
  defparam GSB_CNT_4_3_0_inst.sps_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w10.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w11.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w15.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w16.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w17.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w18.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w20.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w21.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w22.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w23.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w3.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w4.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w5.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w6.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.sps_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.sps_w8.CONF = "01";
  defparam GSB_CNT_4_3_0_inst.sps_w9.CONF = "11";
  defparam GSB_CNT_4_3_0_inst.stub_tbuf3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e0_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e10_w10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e11_w11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e12_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e13_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e14_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e15_w15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e16_w16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e17_w17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e18_w18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e19_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e1_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e20_w20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e21_w21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e22_w22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e23_w23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e2_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e3_w3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e4_w4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e5_w5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e6_w6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e7_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e8_w8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_e9_w9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n0_e20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n0_w5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n10_e6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n10_w15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n11_e11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n11_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n12_e8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n12_w17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n13_e13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n13_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n14_e10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n14_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n15_e15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n15_w16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n16_e12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n16_w21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n17_e17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n17_w18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n18_e14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n18_w23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n19_e19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n19_w20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n1_e1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n1_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n20_e16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n20_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n21_e21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n21_w22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n22_e18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n22_w3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n23_e23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n23_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n2_e22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n2_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n3_e3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n3_w4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n4_e0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n4_w9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n5_e5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n5_w6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n6_e2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n6_w11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n7_e7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n7_w8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n8_e4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n8_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n9_e9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_n9_w10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s0_e22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s0_n0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s0_w2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s10_e4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s10_n10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s10_w8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s11_e9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s11_n11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s11_w13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s12_e10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s12_n12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s12_w14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s13_e15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s13_n13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s13_w19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s14_e8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s14_n14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s14_w12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s15_e13.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s15_n15.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s15_w17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s16_e14.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s16_n16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s16_w18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s17_e19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s17_n17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s17_w23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s18_e12.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s18_n18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s18_w16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s19_e17.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s19_n19.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s19_w21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s1_e3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s1_n1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s1_w7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s20_e18.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s20_n20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s20_w22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s21_e23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s21_n21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s21_w3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s22_e16.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s22_n22.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s22_w20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s23_e21.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s23_n23.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s23_w1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s2_e20.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s2_n2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s2_w0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s3_e1.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s3_n3.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s3_w5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s4_e2.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s4_n4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s4_w6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s5_e7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s5_n5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s5_w11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s6_e0.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s6_n6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s6_w4.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s7_e5.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s7_n7.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s7_w9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s8_e6.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s8_n8.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s8_w10.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s9_e11.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s9_n9.CONF = "1";
  defparam GSB_CNT_4_3_0_inst.switch_s9_w15.CONF = "1";
  GSB_CNT GSB_CNT_4_3_0_inst (
    .E0(),
    .E1(),
    .E2(),
    .E3(),
    .E4(),
    .E5(),
    .E6(),
    .E7(),
    .E8(),
    .E9(),
    .E10(),
    .E11(),
    .E12(),
    .E13(),
    .E14(),
    .E15(),
    .E16(),
    .E17(),
    .E18(),
    .E19(),
    .E20(),
    .E21(),
    .E22(),
    .E23(),
    .N0(),
    .N1(),
    .N2(),
    .N3(),
    .N4(),
    .N5(),
    .N6(),
    .N7(),
    .N8(),
    .N9(),
    .N10(),
    .N11(),
    .N12(),
    .N13(),
    .N14(),
    .N15(),
    .N16(),
    .N17(),
    .N18(),
    .N19(),
    .N20(),
    .N21(),
    .N22(),
    .N23(),
    .W0(),
    .W1(),
    .W2(),
    .W3(),
    .W4(),
    .W5(),
    .W6(),
    .W7(),
    .W8(\net_lcd_db_reg[0]_W8_to_LEFT_E84_2_0 ),
    .W9(),
    .W10(),
    .W11(),
    .W12(),
    .W13(),
    .W14(),
    .W15(),
    .W16(),
    .W17(),
    .W18(),
    .W19(),
    .W20(),
    .W21(),
    .W22(),
    .W23(),
    .S0(),
    .S1(),
    .S2(),
    .S3(),
    .S4(),
    .S5(),
    .S6(),
    .S7(),
    .S8(),
    .S9(),
    .S10(),
    .S11(),
    .S12(),
    .S13(),
    .S14(),
    .S15(),
    .S16(),
    .S17(),
    .S18(),
    .S19(),
    .S20(),
    .S21(),
    .S22(),
    .S23(),
    .H6E0(),
    .H6E1(),
    .H6E2(),
    .H6E3(),
    .H6E4(),
    .H6E5(),
    .H6E6(),
    .H6E7(),
    .H6E8(),
    .H6E9(),
    .H6E10(),
    .H6E11(),
    .H6M0(),
    .H6M1(),
    .H6M2(),
    .H6M3(),
    .H6M4(),
    .H6M5(),
    .H6M6(),
    .H6M7(),
    .H6M8(),
    .H6M9(),
    .H6M10(),
    .H6M11(),
    .H6W0(),
    .H6W1(),
    .H6W2(),
    .H6W3(),
    .H6W4(),
    .H6W5(),
    .H6W6(),
    .H6W7(),
    .H6W8(),
    .H6W9(),
    .H6W10(),
    .H6W11(),
    .LLH0(),
    .LLH6(),
    .GCLK3(),
    .GCLK2(),
    .GCLK1(),
    .GCLK0(),
    .OUT0(),
    .OUT1(),
    .OUT6(),
    .OUT7(),
    .OUT_W0(),
    .OUT_W1(),
    .OUT_E6(),
    .OUT_E7(),
    .TBUF0(),
    .TBUF1(),
    .TBUF2(),
    .TBUF3(),
    .TBUF_STUB3(),
    .V6N0(),
    .V6N1(),
    .V6N2(),
    .V6N3(),
    .V6N4(),
    .V6N5(),
    .V6N6(),
    .V6N7(),
    .V6N8(),
    .V6N9(),
    .V6N10(),
    .V6N11(),
    .V6M0(),
    .V6M1(\net_lcd_db_reg[0]_V6N1_to_V6M14_3_0 ),
    .V6M2(),
    .V6M3(),
    .V6M4(),
    .V6M5(),
    .V6M6(),
    .V6M7(),
    .V6M8(),
    .V6M9(),
    .V6M10(),
    .V6M11(),
    .V6S0(),
    .V6S1(),
    .V6S2(),
    .V6S3(),
    .V6S4(),
    .V6S5(),
    .V6S6(),
    .V6S7(),
    .V6S8(),
    .V6S9(),
    .V6S10(),
    .V6S11(),
    .V6A0(),
    .V6A1(),
    .V6A2(),
    .V6A3(),
    .V6B0(),
    .V6B1(),
    .V6B2(),
    .V6B3(),
    .V6C0(),
    .V6C1(),
    .V6C2(),
    .V6C3(),
    .V6D0(),
    .V6D1(),
    .V6D2(),
    .V6D3(),
    .LLV0(),
    .LLV6(),
    .S0_F_B1(),
    .S0_F_B2(),
    .S0_F_B3(),
    .S0_F_B4(),
    .S0_G_B1(),
    .S0_G_B2(),
    .S0_G_B3(),
    .S0_G_B4(),
    .S0_BX_B(),
    .S0_BY_B(),
    .S0_CE_B(),
    .S0_CLK_B(),
    .S0_SR_B(),
    .S0_X(),
    .S0_XB(),
    .S0_Y(),
    .S0_YB(),
    .S0_XQ(),
    .S0_YQ(),
    .CO_0_LOCAL(),
    .CO_0(),
    .S0_F5(),
    .S0_F5IN(),
    .S1_F_B1(),
    .S1_F_B2(),
    .S1_F_B3(),
    .S1_F_B4(),
    .S1_G_B1(),
    .S1_G_B2(),
    .S1_G_B3(),
    .S1_G_B4(),
    .S1_BX_B(),
    .S1_BY_B(),
    .S1_CE_B(),
    .S1_CLK_B(),
    .S1_SR_B(),
    .S1_X(),
    .S1_XB(),
    .S1_Y(),
    .S1_YB(),
    .S1_XQ(),
    .S1_YQ(),
    .TS_B0(),
    .TS_B1(),
    .CO_1_LOCAL(),
    .CO_1(),
    .S1_F5(),
    .S1_F5IN(),
    .TBUF_OUT0(),
    .TBUF_OUT1(),
    .T_IN0(),
    .T_IN1(),
    .CIN_0_I(),
    .CIN_0_O(),
    .CIN_1_I(),
    .CIN_1_O()
  );

  defparam GSB_LFT_4_2_0_inst.sps_e0.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e1.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e10.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e11.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e12.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e13.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e14.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e15.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e16.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e17.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e18.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e19.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e2.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e20.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e21.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e22.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e23.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e3.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e4.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e5.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e6.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_e7.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e8.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_e9.CONF = "111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e0.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e11.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e5.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e7.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6e9.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_llh0.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh6.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llv0.CONF = "1111111111";
  defparam GSB_LFT_4_2_0_inst.sps_llv6.CONF = "1111111111";
  defparam GSB_LFT_4_2_0_inst.sps_out0.CONF = "1111";
  defparam GSB_LFT_4_2_0_inst.sps_out1.CONF = "1111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n0.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n1.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n2.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6n3.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s0.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s1.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s2.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_v6s3.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.spbu_tbufo0.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.spbu_tbufo1.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.spbu_tbufo2.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.spbu_tbufo3.CONF = "1";
  defparam GSB_LFT_4_2_0_inst.sps_clk1.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_clk2.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_clk3.CONF = "11111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a11.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a5.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a7.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6a9.CONF = "111111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6b3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6c3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6d3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m0.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m1.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m2.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_h6m3.CONF = "11111";
  defparam GSB_LFT_4_2_0_inst.sps_ice1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ice2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ice3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_llh1.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh10.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh11.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh2.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh3.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh4.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh5.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh7.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh8.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_llh9.CONF = "11";
  defparam GSB_LFT_4_2_0_inst.sps_o1.CONF = "110000111";
  defparam GSB_LFT_4_2_0_inst.sps_o2.CONF = "111111111";
  defparam GSB_LFT_4_2_0_inst.sps_o3.CONF = "111111111";
  defparam GSB_LFT_4_2_0_inst.sps_oce1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_oce2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_oce3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_sr_b1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_sr_b2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_sr_b3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_t1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_t2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_t3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_tce1.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_tce2.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_tce3.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ti0_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ti1_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ts0_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.sps_ts1_b.CONF = "1111111";
  defparam GSB_LFT_4_2_0_inst.stub_tbuf1.CONF = "1";
  GSB_LFT GSB_LFT_4_2_0_inst (
    .LEFT_E23(),
    .LEFT_E22(),
    .LEFT_E21(),
    .LEFT_E20(),
    .LEFT_E19(),
    .LEFT_E18(),
    .LEFT_E17(),
    .LEFT_E16(),
    .LEFT_E15(),
    .LEFT_E14(),
    .LEFT_E13(),
    .LEFT_E12(),
    .LEFT_E11(),
    .LEFT_E10(),
    .LEFT_E9(),
    .LEFT_E8(\net_lcd_db_reg[0]_W8_to_LEFT_E84_2_0 ),
    .LEFT_E7(),
    .LEFT_E6(),
    .LEFT_E5(),
    .LEFT_E4(),
    .LEFT_E3(),
    .LEFT_E2(),
    .LEFT_E1(),
    .LEFT_E0(),
    .LEFT_H6E0(),
    .LEFT_H6E1(),
    .LEFT_H6E2(),
    .LEFT_H6E3(),
    .LEFT_H6E4(),
    .LEFT_H6E5(),
    .LEFT_H6E6(),
    .LEFT_H6E7(),
    .LEFT_H6E8(),
    .LEFT_H6E9(),
    .LEFT_H6E10(),
    .LEFT_H6E11(),
    .LEFT_H6A0(),
    .LEFT_H6A1(),
    .LEFT_H6A2(),
    .LEFT_H6A3(),
    .LEFT_H6A4(),
    .LEFT_H6A5(),
    .LEFT_H6A6(),
    .LEFT_H6A7(),
    .LEFT_H6A8(),
    .LEFT_H6A9(),
    .LEFT_H6A10(),
    .LEFT_H6A11(),
    .LEFT_H6B0(),
    .LEFT_H6B1(),
    .LEFT_H6B2(),
    .LEFT_H6B3(),
    .LEFT_H6B4(),
    .LEFT_H6B5(),
    .LEFT_H6B6(),
    .LEFT_H6B7(),
    .LEFT_H6B8(),
    .LEFT_H6B9(),
    .LEFT_H6B10(),
    .LEFT_H6B11(),
    .LEFT_H6M0(),
    .LEFT_H6M1(),
    .LEFT_H6M2(),
    .LEFT_H6M3(),
    .LEFT_H6M4(),
    .LEFT_H6M5(),
    .LEFT_H6M6(),
    .LEFT_H6M7(),
    .LEFT_H6M8(),
    .LEFT_H6M9(),
    .LEFT_H6M10(),
    .LEFT_H6M11(),
    .LEFT_H6C0(),
    .LEFT_H6C1(),
    .LEFT_H6C2(),
    .LEFT_H6C3(),
    .LEFT_H6C4(),
    .LEFT_H6C5(),
    .LEFT_H6C6(),
    .LEFT_H6C7(),
    .LEFT_H6C8(),
    .LEFT_H6C9(),
    .LEFT_H6C10(),
    .LEFT_H6C11(),
    .LEFT_H6D0(),
    .LEFT_H6D1(),
    .LEFT_H6D2(),
    .LEFT_H6D3(),
    .LEFT_H6D4(),
    .LEFT_H6D5(),
    .LEFT_H6D6(),
    .LEFT_H6D7(),
    .LEFT_H6D8(),
    .LEFT_H6D9(),
    .LEFT_H6D10(),
    .LEFT_H6D11(),
    .LEFT_LLH0(),
    .LEFT_LLH1(),
    .LEFT_LLH2(),
    .LEFT_LLH3(),
    .LEFT_LLH4(),
    .LEFT_LLH5(),
    .LEFT_LLH6(),
    .LEFT_LLH7(),
    .LEFT_LLH8(),
    .LEFT_LLH9(),
    .LEFT_LLH10(),
    .LEFT_LLH11(),
    .LEFT_GCLK0(),
    .LEFT_GCLK1(),
    .LEFT_GCLK2(),
    .LEFT_GCLK3(),
    .LEFT_OUT0(),
    .LEFT_OUT1(),
    .LEFT_OUT_E6(),
    .LEFT_OUT_E7(),
    .LEFT_TBUF1_STUB(),
    .LEFT_TBUFO2(),
    .LEFT_TBUFO3(),
    .LEFT_TBUFO0(),
    .LEFT_V6N0(),
    .LEFT_V6N1(),
    .LEFT_V6N2(),
    .LEFT_V6N3(),
    .LEFT_V6A0(),
    .LEFT_V6A1(),
    .LEFT_V6A2(),
    .LEFT_V6A3(),
    .LEFT_V6B0(),
    .LEFT_V6B1(),
    .LEFT_V6B2(),
    .LEFT_V6B3(),
    .LEFT_V6M0(),
    .LEFT_V6M1(),
    .LEFT_V6M2(),
    .LEFT_V6M3(),
    .LEFT_V6C0(),
    .LEFT_V6C1(),
    .LEFT_V6C2(),
    .LEFT_V6C3(),
    .LEFT_V6D0(),
    .LEFT_V6D1(),
    .LEFT_V6D2(),
    .LEFT_V6D3(),
    .LEFT_V6S0(),
    .LEFT_V6S1(),
    .LEFT_V6S2(),
    .LEFT_V6S3(),
    .LEFT_LLV0(),
    .LEFT_LLV6(),
    .LEFT_PCI_CE(),
    .LEFT_I1(),
    .LEFT_I2(),
    .LEFT_I3(),
    .LEFT_IQ1(),
    .LEFT_IQ2(),
    .LEFT_IQ3(),
    .LEFT_ICE1(),
    .LEFT_ICE2(),
    .LEFT_ICE3(),
    .LEFT_O1(\net_lcd_db_reg[0]_LEFT_O1_to_OUT4_2_0 ),
    .LEFT_O2(),
    .LEFT_O3(),
    .LEFT_OCE1(),
    .LEFT_OCE2(),
    .LEFT_OCE3(),
    .LEFT_T1(),
    .LEFT_T2(),
    .LEFT_T3(),
    .LEFT_TCE1(),
    .LEFT_TCE2(),
    .LEFT_TCE3(),
    .LEFT_CLK1(),
    .LEFT_CLK2(),
    .LEFT_CLK3(),
    .LEFT_SR_B1(),
    .LEFT_SR_B2(),
    .LEFT_SR_B3(),
    .LEFT_TS0_B(),
    .LEFT_TS1_B(),
    .LEFT_TO0(),
    .LEFT_TO1(),
    .LEFT_TI0_B(),
    .LEFT_TI1_B()
  );

  GSB_CLKC GSB_CLKC_18_28_0_inst (
    .CLKC_GCLK0(),
    .CLKC_GCLK1(\net_IBuf-clkpad-clk_CLKB_GCLK1_to_CLKC_GCLK118_28_0 ),
    .CLKC_GCLK2(),
    .CLKC_GCLK3(),
    .CLKC_HGCLK0(),
    .CLKC_HGCLK1(\net_IBuf-clkpad-clk_CLKC_HGCLK1_to_BRAM_CLKH_GCLK118_1_0 ),
    .CLKC_HGCLK2(),
    .CLKC_HGCLK3(),
    .CLKC_VGCLK0(),
    .CLKC_VGCLK1(),
    .CLKC_VGCLK2(),
    .CLKC_VGCLK3()
  );

  GSB_CLKL GSB_CLKL_18_1_0_inst (
    .BRAM_CLKH_GCLK0(),
    .BRAM_CLKH_GCLK1(\net_IBuf-clkpad-clk_CLKC_HGCLK1_to_BRAM_CLKH_GCLK118_1_0 ),
    .BRAM_CLKH_GCLK2(),
    .BRAM_CLKH_GCLK3(),
    .BRAM_CLKH_VGCLK0(),
    .BRAM_CLKH_VGCLK1(\net_IBuf-clkpad-clk_BRAM_CLKH_VGCLK1_to_BRAM_GCLKIN17_1_0 ),
    .BRAM_CLKH_VGCLK2(),
    .BRAM_CLKH_VGCLK3()
  );

  defparam GSB_LBRAMB_7_1_0_inst.sps_llv6.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.spbu_gclk_clbb0.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.spbu_gclk_clbb1.CONF = "0";
  defparam GSB_LBRAMB_7_1_0_inst.spbu_gclk_clbb2.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.spbu_gclk_clbb3.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.spbu_gclk_iobb0.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.spbu_gclk_iobb1.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.spbu_gclk_iobb2.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.spbu_gclk_iobb3.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.sps_addra0.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_addra1.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_addra2.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_addra3.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_addrb0.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_addrb1.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_addrb2.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_addrb3.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_clka.CONF = "1111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_dia1.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_dia11.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_dia3.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_dia9.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_dib1.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_dib11.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_dib3.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_dib9.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb0.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb1.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb10.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb11.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb12.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb13.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb14.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb15.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb16.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb17.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb18.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb19.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb2.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb20.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb21.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb22.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb23.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb3.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb4.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb5.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb6.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb7.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb8.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_eb9.CONF = "11";
  defparam GSB_LBRAMB_7_1_0_inst.sps_h6bb0.CONF = "111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_h6bb1.CONF = "111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_h6bb2.CONF = "111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_h6bb3.CONF = "111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_h6mb0.CONF = "111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_h6mb1.CONF = "111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_h6mb2.CONF = "111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_h6mb3.CONF = "111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_lhb0.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_lhb3.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_lhb6.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_lhb9.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_llv10.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_llv2.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_raddrs10.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_raddrs14.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_raddrs18.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_raddrs2.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_raddrs22.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_raddrs26.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_raddrs30.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_raddrs6.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_rdins10.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_rdins14.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_rdins18.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_rdins2.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_rdins22.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_rdins26.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_rdins30.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_rdins6.CONF = "111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_rsta.CONF = "1111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_sela.CONF = "1111111";
  defparam GSB_LBRAMB_7_1_0_inst.sps_wea.CONF = "1111111";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa13_rdouts0.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa13_rdouts17.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa1_rdouts23.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa1_rdouts24.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa1_rdouts5.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa1_rdouts6.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa5_rdouts0.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa5_rdouts15.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa5_rdouts17.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa5_rdouts18.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa9_rdouts23.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_doa9_rdouts6.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob13_rdouts1.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob13_rdouts18.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob1_rdouts24.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob1_rdouts25.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob1_rdouts6.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob1_rdouts7.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob5_rdouts0.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob5_rdouts1.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob5_rdouts18.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob5_rdouts19.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob9_rdouts24.CONF = "1";
  defparam GSB_LBRAMB_7_1_0_inst.tribuf_dob9_rdouts7.CONF = "1";
  GSB_LBRAMB GSB_LBRAMB_7_1_0_inst (
    .BRAM_EB0(),
    .BRAM_EB1(),
    .BRAM_EB2(),
    .BRAM_EB3(),
    .BRAM_EB4(),
    .BRAM_EB5(),
    .BRAM_EB6(),
    .BRAM_EB7(),
    .BRAM_EB8(),
    .BRAM_EB9(),
    .BRAM_EB10(),
    .BRAM_EB11(),
    .BRAM_EB12(),
    .BRAM_EB13(),
    .BRAM_EB14(),
    .BRAM_EB15(),
    .BRAM_EB16(),
    .BRAM_EB17(),
    .BRAM_EB18(),
    .BRAM_EB19(),
    .BRAM_EB20(),
    .BRAM_EB21(),
    .BRAM_EB22(),
    .BRAM_EB23(),
    .BRAM_H6EB0(),
    .BRAM_H6EB1(),
    .BRAM_H6EB2(),
    .BRAM_H6EB3(),
    .BRAM_H6BB0(),
    .BRAM_H6BB1(),
    .BRAM_H6BB2(),
    .BRAM_H6BB3(),
    .BRAM_H6MB0(),
    .BRAM_H6MB1(),
    .BRAM_H6MB2(),
    .BRAM_H6MB3(),
    .BRAM_H6DB0(),
    .BRAM_H6DB1(),
    .BRAM_H6DB2(),
    .BRAM_H6DB3(),
    .BRAM_LHB0(),
    .BRAM_LHB3(),
    .BRAM_LHB6(),
    .BRAM_LHB9(),
    .BRAM_LLV0(),
    .BRAM_LLV1(),
    .BRAM_LLV2(),
    .BRAM_LLV3(),
    .BRAM_LLV4(),
    .BRAM_LLV5(),
    .BRAM_LLV6(),
    .BRAM_LLV7(),
    .BRAM_LLV8(),
    .BRAM_LLV9(),
    .BRAM_LLV10(),
    .BRAM_LLV11(),
    .BRAM_GCLKIN0(),
    .BRAM_GCLKIN1(\net_IBuf-clkpad-clk_BRAM_CLKH_VGCLK1_to_BRAM_GCLKIN17_1_0 ),
    .BRAM_GCLKIN2(),
    .BRAM_GCLKIN3(),
    .BRAM_GCLK_IOBB0(),
    .BRAM_GCLK_IOBB1(),
    .BRAM_GCLK_IOBB2(),
    .BRAM_GCLK_IOBB3(),
    .BRAM_GCLK_CLBB0(),
    .BRAM_GCLK_CLBB1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBB1_to_GCLK17_3_0 ),
    .BRAM_GCLK_CLBB2(),
    .BRAM_GCLK_CLBB3(),
    .BRAM_RDOUTS0(),
    .BRAM_RDOUTS1(),
    .BRAM_RDOUTS2(),
    .BRAM_RDOUTS5(),
    .BRAM_RDOUTS6(),
    .BRAM_RDOUTS7(),
    .BRAM_RDOUTS10(),
    .BRAM_RDOUTS14(),
    .BRAM_RDOUTS15(),
    .BRAM_RDOUTS17(),
    .BRAM_RDOUTS18(),
    .BRAM_RDOUTS19(),
    .BRAM_RDOUTS22(),
    .BRAM_RDOUTS23(),
    .BRAM_RDOUTS24(),
    .BRAM_RDOUTS25(),
    .BRAM_RDOUTS26(),
    .BRAM_RDOUTS30(),
    .BRAM_RDINS2(),
    .BRAM_RDINS6(),
    .BRAM_RDINS7(),
    .BRAM_RDINS8(),
    .BRAM_RDINS9(),
    .BRAM_RDINS10(),
    .BRAM_RDINS11(),
    .BRAM_RDINS12(),
    .BRAM_RDINS13(),
    .BRAM_RDINS14(),
    .BRAM_RDINS18(),
    .BRAM_RDINS22(),
    .BRAM_RDINS25(),
    .BRAM_RDINS26(),
    .BRAM_RDINS27(),
    .BRAM_RDINS29(),
    .BRAM_RDINS30(),
    .BRAM_RDINS31(),
    .BRAM_RADDRS0(),
    .BRAM_RADDRS1(),
    .BRAM_RADDRS2(),
    .BRAM_RADDRS3(),
    .BRAM_RADDRS4(),
    .BRAM_RADDRS5(),
    .BRAM_RADDRS6(),
    .BRAM_RADDRS7(),
    .BRAM_RADDRS8(),
    .BRAM_RADDRS9(),
    .BRAM_RADDRS10(),
    .BRAM_RADDRS11(),
    .BRAM_RADDRS14(),
    .BRAM_RADDRS18(),
    .BRAM_RADDRS22(),
    .BRAM_RADDRS24(),
    .BRAM_RADDRS25(),
    .BRAM_RADDRS26(),
    .BRAM_RADDRS27(),
    .BRAM_RADDRS28(),
    .BRAM_RADDRS29(),
    .BRAM_RADDRS30(),
    .BRAM_RADDRS31(),
    .BRAM_DIA1(),
    .BRAM_DIA3(),
    .BRAM_DIA9(),
    .BRAM_DIA11(),
    .BRAM_DIB1(),
    .BRAM_DIB3(),
    .BRAM_DIB9(),
    .BRAM_DIB11(),
    .BRAM_DOA1(),
    .BRAM_DOA5(),
    .BRAM_DOA9(),
    .BRAM_DOA13(),
    .BRAM_DOB1(),
    .BRAM_DOB5(),
    .BRAM_DOB9(),
    .BRAM_DOB13(),
    .BRAM_ADDRA0(),
    .BRAM_ADDRA1(),
    .BRAM_ADDRA2(),
    .BRAM_ADDRA3(),
    .BRAM_ADDRB0(),
    .BRAM_ADDRB1(),
    .BRAM_ADDRB2(),
    .BRAM_ADDRB3(),
    .BRAM_CLKA(),
    .BRAM_WEA(),
    .BRAM_SELA(),
    .BRAM_RSTA()
  );

  defparam GSB_LBRAMD_9_1_0_inst.sps_llv0.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.spbu_gclk_clbd0.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.spbu_gclk_clbd1.CONF = "0";
  defparam GSB_LBRAMD_9_1_0_inst.spbu_gclk_clbd2.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.spbu_gclk_clbd3.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.spbu_gclk_iobd0.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.spbu_gclk_iobd1.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.spbu_gclk_iobd2.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.spbu_gclk_iobd3.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.sps_addra10.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_addra11.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_addra8.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_addra9.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_addrb10.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_addrb11.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_addrb8.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_addrb9.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_dia14.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_dia15.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_dia6.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_dia7.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_dib14.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_dib15.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_dib6.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_dib7.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed0.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed1.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed10.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed11.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed12.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed13.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed14.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed15.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed16.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed17.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed18.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed19.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed2.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed20.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed21.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed22.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed23.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed3.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed4.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed5.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed6.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed7.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed8.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_ed9.CONF = "11";
  defparam GSB_LBRAMD_9_1_0_inst.sps_h6bd0.CONF = "111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_h6bd1.CONF = "111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_h6bd2.CONF = "111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_h6bd3.CONF = "111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_h6md0.CONF = "111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_h6md1.CONF = "111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_h6md2.CONF = "111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_h6md3.CONF = "111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_lhd0.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_lhd3.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_lhd6.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_lhd9.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_llv4.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_llv8.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_raddrs0.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_raddrs12.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_raddrs16.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_raddrs20.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_raddrs24.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_raddrs28.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_raddrs4.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_raddrs8.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_rdins0.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_rdins12.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_rdins16.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_rdins20.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_rdins24.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_rdins28.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_rdins4.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.sps_rdins8.CONF = "111111";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa11_rdouts19.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa11_rdouts2.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa15_rdouts25.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa15_rdouts8.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa3_rdouts1.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa3_rdouts19.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa3_rdouts2.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa3_rdouts20.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa7_rdouts25.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa7_rdouts26.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa7_rdouts7.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_doa7_rdouts8.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob11_rdouts20.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob11_rdouts3.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob15_rdouts26.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob15_rdouts9.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob3_rdouts2.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob3_rdouts20.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob3_rdouts21.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob3_rdouts3.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob7_rdouts26.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob7_rdouts27.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob7_rdouts8.CONF = "1";
  defparam GSB_LBRAMD_9_1_0_inst.tribuf_dob7_rdouts9.CONF = "1";
  GSB_LBRAMD GSB_LBRAMD_9_1_0_inst (
    .BRAM_ED0(),
    .BRAM_ED1(),
    .BRAM_ED2(),
    .BRAM_ED3(),
    .BRAM_ED4(),
    .BRAM_ED5(),
    .BRAM_ED6(),
    .BRAM_ED7(),
    .BRAM_ED8(),
    .BRAM_ED9(),
    .BRAM_ED10(),
    .BRAM_ED11(),
    .BRAM_ED12(),
    .BRAM_ED13(),
    .BRAM_ED14(),
    .BRAM_ED15(),
    .BRAM_ED16(),
    .BRAM_ED17(),
    .BRAM_ED18(),
    .BRAM_ED19(),
    .BRAM_ED20(),
    .BRAM_ED21(),
    .BRAM_ED22(),
    .BRAM_ED23(),
    .BRAM_H6ED0(),
    .BRAM_H6ED1(),
    .BRAM_H6ED2(),
    .BRAM_H6ED3(),
    .BRAM_H6BD0(),
    .BRAM_H6BD1(),
    .BRAM_H6BD2(),
    .BRAM_H6BD3(),
    .BRAM_H6MD0(),
    .BRAM_H6MD1(),
    .BRAM_H6MD2(),
    .BRAM_H6MD3(),
    .BRAM_H6DD0(),
    .BRAM_H6DD1(),
    .BRAM_H6DD2(),
    .BRAM_H6DD3(),
    .BRAM_LHD0(),
    .BRAM_LHD3(),
    .BRAM_LHD6(),
    .BRAM_LHD9(),
    .BRAM_LLV0(),
    .BRAM_LLV4(),
    .BRAM_LLV8(),
    .BRAM_RDOUTS0(),
    .BRAM_RDOUTS1(),
    .BRAM_RDOUTS2(),
    .BRAM_RDOUTS3(),
    .BRAM_RDOUTS4(),
    .BRAM_RDOUTS7(),
    .BRAM_RDOUTS8(),
    .BRAM_RDOUTS9(),
    .BRAM_RDOUTS12(),
    .BRAM_RDOUTS16(),
    .BRAM_RDOUTS19(),
    .BRAM_RDOUTS20(),
    .BRAM_RDOUTS21(),
    .BRAM_RDOUTS24(),
    .BRAM_RDOUTS25(),
    .BRAM_RDOUTS26(),
    .BRAM_RDOUTS27(),
    .BRAM_RDOUTS28(),
    .BRAM_RADDRS0(),
    .BRAM_RADDRS4(),
    .BRAM_RADDRS8(),
    .BRAM_RADDRS12(),
    .BRAM_RADDRS16(),
    .BRAM_RADDRS17(),
    .BRAM_RADDRS18(),
    .BRAM_RADDRS19(),
    .BRAM_RADDRS20(),
    .BRAM_RADDRS21(),
    .BRAM_RADDRS22(),
    .BRAM_RADDRS23(),
    .BRAM_RADDRS24(),
    .BRAM_RADDRS25(),
    .BRAM_RADDRS26(),
    .BRAM_RADDRS27(),
    .BRAM_RADDRS28(),
    .BRAM_RDINS0(),
    .BRAM_RDINS4(),
    .BRAM_RDINS8(),
    .BRAM_RDINS9(),
    .BRAM_RDINS10(),
    .BRAM_RDINS11(),
    .BRAM_RDINS12(),
    .BRAM_RDINS13(),
    .BRAM_RDINS14(),
    .BRAM_RDINS15(),
    .BRAM_RDINS16(),
    .BRAM_RDINS17(),
    .BRAM_RDINS20(),
    .BRAM_RDINS24(),
    .BRAM_RDINS27(),
    .BRAM_RDINS28(),
    .BRAM_RDINS29(),
    .BRAM_RDINS31(),
    .BRAM_GCLKIN0(),
    .BRAM_GCLKIN1(\net_IBuf-clkpad-clk_BRAM_CLKH_VGCLK1_to_BRAM_GCLKIN17_1_0 ),
    .BRAM_GCLKIN2(),
    .BRAM_GCLKIN3(),
    .BRAM_GCLK_IOBD0(),
    .BRAM_GCLK_IOBD1(),
    .BRAM_GCLK_IOBD2(),
    .BRAM_GCLK_IOBD3(),
    .BRAM_GCLK_CLBD0(),
    .BRAM_GCLK_CLBD1(\net_IBuf-clkpad-clk_BRAM_GCLK_CLBD1_to_GCLK19_3_0 ),
    .BRAM_GCLK_CLBD2(),
    .BRAM_GCLK_CLBD3(),
    .BRAM_DIA6(),
    .BRAM_DIA7(),
    .BRAM_DIA14(),
    .BRAM_DIA15(),
    .BRAM_DIB6(),
    .BRAM_DIB7(),
    .BRAM_DIB14(),
    .BRAM_DIB15(),
    .BRAM_DOA3(),
    .BRAM_DOA7(),
    .BRAM_DOA11(),
    .BRAM_DOA15(),
    .BRAM_DOB3(),
    .BRAM_DOB7(),
    .BRAM_DOB11(),
    .BRAM_DOB15(),
    .BRAM_ADDRB8(),
    .BRAM_ADDRB9(),
    .BRAM_ADDRB10(),
    .BRAM_ADDRB11(),
    .BRAM_ADDRA8(),
    .BRAM_ADDRA9(),
    .BRAM_ADDRA10(),
    .BRAM_ADDRA11()
  );
endmodule
